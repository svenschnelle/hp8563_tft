library ieee;
use ieee.std_logic_1164.all;
use IEEE.numeric_std.all;

entity charmap is
	port (input: in std_logic_vector(11 downto 0);
	      output: out integer range 0 to 255);
end entity;
architecture rtl of charmap is
begin

output <= 16#20# when input = x"02b" else
	  16#21# when input = x"02c" else
	  16#22# when input = x"032" else
	  16#23# when input = x"037" else
	  16#24# when input = x"044" else
	  16#25# when input = x"052" else
	  16#26# when input = x"05a" else
	  16#27# when input = x"067" else
	  16#28# when input = x"06a" else
	  16#29# when input = x"06f" else
	  16#2a# when input = x"074" else
	  16#2b# when input = x"07b" else
	  16#2c# when input = x"082" else
	  16#2d# when input = x"088" else
	  16#2e# when input = x"08c" else
	  16#2f# when input = x"091" else
	  16#30# when input = x"095" else
	  16#31# when input = x"0a1" else
	  16#32# when input = x"0a8" else
	  16#33# when input = x"0b2" else
	  16#34# when input = x"0be" else
	  16#35# when input = x"0c6" else
	  16#36# when input = x"0d1" else
	  16#37# when input = x"0dc" else
	  16#38# when input = x"0e2" else
	  16#39# when input = x"0ef" else
	  16#3a# when input = x"0fa" else
	  16#3b# when input = x"103" else
	  16#3c# when input = x"10d" else
	  16#3d# when input = x"113" else
	  16#3e# when input = x"11a" else
	  16#3f# when input = x"120" else
	  16#40# when input = x"129" else
	  16#41# when input = x"137" else
	  16#42# when input = x"140" else
	  16#43# when input = x"14e" else
	  16#44# when input = x"157" else
	  16#45# when input = x"160" else
	  16#46# when input = x"16b" else
	  16#47# when input = x"174" else
	  16#48# when input = x"17f" else
	  16#49# when input = x"189" else
	  16#4a# when input = x"191" else
	  16#4b# when input = x"198" else
	  16#4c# when input = x"1a2" else
	  16#4d# when input = x"1a8" else
	  16#4e# when input = x"1b2" else
	  16#4f# when input = x"1ba" else
	  16#50# when input = x"1c5" else
	  16#51# when input = x"1cd" else
	  16#52# when input = x"1da" else
	  16#53# when input = x"1e5" else
	  16#54# when input = x"1ef" else
	  16#55# when input = x"1f6" else
	  16#56# when input = x"1fe" else
	  16#57# when input = x"204" else
	  16#58# when input = x"20e" else
	  16#59# when input = x"215" else
	  16#5a# when input = x"21d" else
	  16#5b# when input = x"225" else
	  16#5c# when input = x"22c" else
	  16#5d# when input = x"230" else
	  16#5e# when input = x"237" else
	  16#5f# when input = x"23d" else
	  16#60# when input = x"241" else
	  16#61# when input = x"244" else
	  16#62# when input = x"24e" else
	  16#63# when input = x"258" else
	  16#64# when input = x"25f" else
	  16#65# when input = x"269" else
	  16#66# when input = x"272" else
	  16#67# when input = x"27a" else
	  16#68# when input = x"286" else
	  16#69# when input = x"28e" else
	  16#6a# when input = x"294" else
	  16#6b# when input = x"29c" else
	  16#6c# when input = x"2a4" else
	  16#6d# when input = x"2a8" else
	  16#6e# when input = x"2b3" else
	  16#6f# when input = x"2ba" else
	  16#70# when input = x"2c2" else
	  16#71# when input = x"2cc" else
	  16#72# when input = x"2d6" else
	  16#73# when input = x"2dc" else
	  16#74# when input = x"2e5" else
	  16#75# when input = x"2ec" else
	  16#76# when input = x"2f3" else
	  16#77# when input = x"2f7" else
	  16#78# when input = x"2fd" else
	  16#79# when input = x"304" else
	  16#7a# when input = x"30c" else
	  16#7b# when input = x"314" else
	  16#7c# when input = x"31c" else
	  16#7d# when input = x"320" else
	  16#7e# when input = x"328" else
	  16#7f# when input = x"399" else
	  16#80# when input = x"32e" else
	  16#81# when input = x"32f" else
	  16#82# when input = x"330" else
	  16#83# when input = x"331" else
	  16#84# when input = x"332" else
	  16#85# when input = x"333" else
	  16#86# when input = x"334" else
	  16#87# when input = x"335" else
	  16#88# when input = x"336" else
	  16#89# when input = x"337" else
	  16#8a# when input = x"338" else
	  16#8b# when input = x"339" else
	  16#8c# when input = x"33a" else
	  16#8d# when input = x"33b" else
	  16#8e# when input = x"33c" else
	  16#8f# when input = x"33d" else
	  16#90# when input = x"33e" else
	  16#91# when input = x"33f" else
	  16#92# when input = x"341" else
	  16#93# when input = x"343" else
	  16#94# when input = x"345" else
	  16#95# when input = x"347" else
	  16#96# when input = x"348" else
	  16#97# when input = x"349" else
	  16#98# when input = x"34a" else
	  16#99# when input = x"34b" else
	  16#9a# when input = x"34c" else
	  16#9b# when input = x"34d" else
	  16#9c# when input = x"34e" else
	  16#9d# when input = x"34f" else
	  16#9e# when input = x"350" else
	  16#9f# when input = x"351" else
	  16#a0# when input = x"352" else
	  16#a1# when input = x"358" else
	  16#a2# when input = x"35c" else
	  16#a3# when input = x"361" else
	  16#a4# when input = x"36b" else
	  16#a5# when input = x"377" else
	  16#a6# when input = x"381" else
	  16#a7# when input = x"38f" else
	  16#a8# when input = x"392" else
	  16#a9# when input = x"399" else
	  16#aa# when input = x"3a0" else
	  16#ab# when input = x"3af" else
	  16#ac# when input = x"3b9" else
	  16#ad# when input = x"3bf" else
	  16#ae# when input = x"3c3" else
	  16#af# when input = x"3c8" else
	  16#b0# when input = x"3d0" else
	  16#b1# when input = x"3d8" else
	  16#b2# when input = x"3db" else
	  16#b3# when input = x"3e1" else
	  16#b4# when input = x"3e8" else
	  16#b5# when input = x"3ed" else
	  16#b6# when input = x"3f3" else
	  16#b7# when input = x"3fa" else
	  16#b8# when input = x"3ff" else
	  16#b9# when input = x"404" else
	  16#ba# when input = x"40c" else
	  16#bb# when input = x"413" else
	  16#bc# when input = x"41a" else
	  16#bd# when input = x"423" else
	  16#be# when input = x"42d" else
	  16#bf# when input = x"436" else
	  16#c0# when input = x"43a" else
	  16#c1# when input = x"440" else
	  16#c2# when input = x"446" else
	  16#c3# when input = x"44f" else
	  16#c4# when input = x"458" else
	  16#c5# when input = x"460" else
	  16#c6# when input = x"461" else
	  16#c7# when input = x"462" else
	  16#c8# when input = x"46d" else
	  16#c9# when input = x"475" else
	  16#ca# when input = x"47a" else
	  16#cb# when input = x"47b" else
	  16#cc# when input = x"47c" else
	  16#cd# when input = x"480" else
	  16#ce# when input = x"487" else
	  16#cf# when input = x"48e" else
	  16#d0# when input = x"496" else
	  16#d1# when input = x"49f" else
	  16#d2# when input = x"4ab" else
	  16#d3# when input = x"4b1" else
	  16#d4# when input = x"4b8" else
	  16#d5# when input = x"4bd" else
	  16#d6# when input = x"4c7" else
	  16#d7# when input = x"4cb" else
	  16#d8# when input = x"4cc" else
	  16#d9# when input = x"4d3" else
	  16#da# when input = x"4da" else
	  16#db# when input = x"4db" else
	  16#dc# when input = x"4e9" else
	  16#dd# when input = x"4f5" else
	  16#de# when input = x"502" else
	  16#df# when input = x"510" else
	  16#e0# when input = x"512" else
	  16#e1# when input = x"51c" else
	  16#e2# when input = x"526" else
	  16#e3# when input = x"534" else
	  16#e4# when input = x"53b" else
	  16#e5# when input = x"546" else
	  16#e6# when input = x"54f" else
	  16#e7# when input = x"559" else
	  16#e8# when input = x"560" else
	  16#e9# when input = x"567" else
	  16#ea# when input = x"56c" else
	  16#eb# when input = x"577" else
	  16#ec# when input = x"57e" else
	  16#ed# when input = x"585" else
	  16#ee# when input = x"590" else
	  16#ef# when input = x"596" else
	  16#f0# when input = x"59e" else
	  16#f1# when input = x"5a6" else
	  16#f2# when input = x"5b2" else
	  16#f3# when input = x"5bb" else
	  16#f4# when input = x"5c4" else
	  16#f5# when input = x"5cb" else
	  16#f6# when input = x"5d3" else
	  16#f7# when input = x"5e0" else
	  16#f8# when input = x"5ea" else
	  16#f9# when input = x"5f4" else
	  16#fa# when input = x"5fc" else
	  16#fb# when input = x"607" else
	  16#fc# when input = x"614" else
	  16#fd# when input = x"61e" else
	  16#fe# when input = x"62a" else
	  16#ff# when input = x"638" else
	 0;
end;
