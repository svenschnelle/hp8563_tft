library ieee;
use ieee.std_logic_1164.all;

entity testrom is
	port(read_clock_i: in std_logic;
	   read_addr_i: in integer range 0 to 8191;
	   read_data_o: out std_logic_vector(15 downto 0)
);
end testrom;
architecture rtl of testrom is
begin
	process (read_clock_i)
	begin
		if (rising_edge(read_clock_i)) then
			case read_addr_i is
				when 0 => read_data_o <= x"a002";
				when 1 => read_data_o <= x"72c0";
				when 2 => read_data_o <= x"021c";
				when 3 => read_data_o <= x"72d0";
				when 4 => read_data_o <= x"021c";
				when 5 => read_data_o <= x"72c0";
				when 6 => read_data_o <= x"01b8";
				when 7 => read_data_o <= x"72d0";
				when 8 => read_data_o <= x"01b8";
				when 9 => read_data_o <= x"72c0";
			       when 10 => read_data_o <= x"0154";
			       when 11 => read_data_o <= x"72d0";
			       when 12 => read_data_o <= x"0154";
			       when 13 => read_data_o <= x"72c0";
			       when 14 => read_data_o <= x"00f0";
			       when 15 => read_data_o <= x"72d0";
			       when 16 => read_data_o <= x"00f0";
			       when 17 => read_data_o <= x"72c0";
			       when 18 => read_data_o <= x"008c";
			       when 19 => read_data_o <= x"72d0";
			       when 20 => read_data_o <= x"008c";
			       when 21 => read_data_o <= x"72c0";
			       when 22 => read_data_o <= x"0028";
			       when 23 => read_data_o <= x"72d0";
			       when 24 => read_data_o <= x"0028";
			       when 25 => read_data_o <= x"a07a";
			       when 26 => read_data_o <= x"a000";
			       when 27 => read_data_o <= x"a000";
			       when 28 => read_data_o <= x"a000";
			       when 29 => read_data_o <= x"a000";
			       when 30 => read_data_o <= x"a000";
			       when 31 => read_data_o <= x"a000";
			       when 32 => read_data_o <= x"a000";
			       when 33 => read_data_o <= x"a000";
			       when 34 => read_data_o <= x"a000";
			       when 35 => read_data_o <= x"a000";
			       when 36 => read_data_o <= x"a000";
			       when 37 => read_data_o <= x"a000";
			       when 38 => read_data_o <= x"a000";
			       when 39 => read_data_o <= x"a000";
			       when 40 => read_data_o <= x"a000";
			       when 41 => read_data_o <= x"a000";
			       when 42 => read_data_o <= x"a000";
			       when 43 => read_data_o <= x"a000";
			       when 44 => read_data_o <= x"a000";
			       when 45 => read_data_o <= x"a000";
			       when 46 => read_data_o <= x"a000";
			       when 47 => read_data_o <= x"a000";
			       when 48 => read_data_o <= x"a000";
			       when 49 => read_data_o <= x"a000";
			       when 50 => read_data_o <= x"a000";
			       when 51 => read_data_o <= x"a000";
			       when 52 => read_data_o <= x"a000";
			       when 53 => read_data_o <= x"a000";
			       when 54 => read_data_o <= x"a000";
			       when 55 => read_data_o <= x"a000";
			       when 56 => read_data_o <= x"a000";
			       when 57 => read_data_o <= x"a000";
			       when 58 => read_data_o <= x"a000";
			       when 59 => read_data_o <= x"a000";
			       when 60 => read_data_o <= x"a000";
			       when 61 => read_data_o <= x"a0a2";
			       when 62 => read_data_o <= x"0094";
			       when 63 => read_data_o <= x"d02b";
			       when 64 => read_data_o <= x"a000";
			       when 65 => read_data_o <= x"a000";
			       when 66 => read_data_o <= x"a000";
			       when 67 => read_data_o <= x"a000";
			       when 68 => read_data_o <= x"a000";
			       when 69 => read_data_o <= x"a000";
			       when 70 => read_data_o <= x"a000";
			       when 71 => read_data_o <= x"a000";
			       when 72 => read_data_o <= x"a000";
			       when 73 => read_data_o <= x"a000";
			       when 74 => read_data_o <= x"a000";
			       when 75 => read_data_o <= x"a000";
			       when 76 => read_data_o <= x"a000";
			       when 77 => read_data_o <= x"a000";
			       when 78 => read_data_o <= x"a000";
			       when 79 => read_data_o <= x"a000";
			       when 80 => read_data_o <= x"a000";
			       when 81 => read_data_o <= x"a0ca";
			       when 82 => read_data_o <= x"0094";
			       when 83 => read_data_o <= x"d02b";
			       when 84 => read_data_o <= x"a000";
			       when 85 => read_data_o <= x"a000";
			       when 86 => read_data_o <= x"a000";
			       when 87 => read_data_o <= x"a000";
			       when 88 => read_data_o <= x"a000";
			       when 89 => read_data_o <= x"a000";
			       when 90 => read_data_o <= x"a000";
			       when 91 => read_data_o <= x"a000";
			       when 92 => read_data_o <= x"a000";
			       when 93 => read_data_o <= x"a000";
			       when 94 => read_data_o <= x"a000";
			       when 95 => read_data_o <= x"a000";
			       when 96 => read_data_o <= x"a000";
			       when 97 => read_data_o <= x"a000";
			       when 98 => read_data_o <= x"a000";
			       when 99 => read_data_o <= x"a000";
			      when 100 => read_data_o <= x"a000";
			      when 101 => read_data_o <= x"72c0";
			      when 102 => read_data_o <= x"02dc";
			      when 103 => read_data_o <= x"d02b";
			      when 104 => read_data_o <= x"d02b";
			      when 105 => read_data_o <= x"d02b";
			      when 106 => read_data_o <= x"d02b";
			      when 107 => read_data_o <= x"d02b";
			      when 108 => read_data_o <= x"d02b";
			      when 109 => read_data_o <= x"d02b";
			      when 110 => read_data_o <= x"d02b";
			      when 111 => read_data_o <= x"72c0";
			      when 112 => read_data_o <= x"0294";
			      when 113 => read_data_o <= x"d02b";
			      when 114 => read_data_o <= x"d02b";
			      when 115 => read_data_o <= x"d02b";
			      when 116 => read_data_o <= x"d02b";
			      when 117 => read_data_o <= x"d02b";
			      when 118 => read_data_o <= x"d02b";
			      when 119 => read_data_o <= x"d02b";
			      when 120 => read_data_o <= x"d02b";
			      when 121 => read_data_o <= x"72c0";
			      when 122 => read_data_o <= x"027c";
			      when 123 => read_data_o <= x"d02b";
			      when 124 => read_data_o <= x"d02b";
			      when 125 => read_data_o <= x"d02b";
			      when 126 => read_data_o <= x"d02b";
			      when 127 => read_data_o <= x"d02b";
			      when 128 => read_data_o <= x"d02b";
			      when 129 => read_data_o <= x"d02b";
			      when 130 => read_data_o <= x"d02b";
			      when 131 => read_data_o <= x"72c0";
			      when 132 => read_data_o <= x"0230";
			      when 133 => read_data_o <= x"d02b";
			      when 134 => read_data_o <= x"d02b";
			      when 135 => read_data_o <= x"d02b";
			      when 136 => read_data_o <= x"d02b";
			      when 137 => read_data_o <= x"d02b";
			      when 138 => read_data_o <= x"d02b";
			      when 139 => read_data_o <= x"d02b";
			      when 140 => read_data_o <= x"d02b";
			      when 141 => read_data_o <= x"72c0";
			      when 142 => read_data_o <= x"0218";
			      when 143 => read_data_o <= x"d02b";
			      when 144 => read_data_o <= x"d02b";
			      when 145 => read_data_o <= x"d02b";
			      when 146 => read_data_o <= x"d02b";
			      when 147 => read_data_o <= x"d02b";
			      when 148 => read_data_o <= x"d02b";
			      when 149 => read_data_o <= x"d02b";
			      when 150 => read_data_o <= x"d02b";
			      when 151 => read_data_o <= x"72c0";
			      when 152 => read_data_o <= x"01cc";
			      when 153 => read_data_o <= x"d02b";
			      when 154 => read_data_o <= x"d02b";
			      when 155 => read_data_o <= x"d02b";
			      when 156 => read_data_o <= x"d02b";
			      when 157 => read_data_o <= x"d02b";
			      when 158 => read_data_o <= x"d02b";
			      when 159 => read_data_o <= x"d02b";
			      when 160 => read_data_o <= x"d02b";
			      when 161 => read_data_o <= x"72c0";
			      when 162 => read_data_o <= x"01b4";
			      when 163 => read_data_o <= x"d02b";
			      when 164 => read_data_o <= x"d02b";
			      when 165 => read_data_o <= x"d02b";
			      when 166 => read_data_o <= x"d02b";
			      when 167 => read_data_o <= x"d02b";
			      when 168 => read_data_o <= x"d02b";
			      when 169 => read_data_o <= x"d02b";
			      when 170 => read_data_o <= x"d02b";
			      when 171 => read_data_o <= x"72c0";
			      when 172 => read_data_o <= x"0168";
			      when 173 => read_data_o <= x"d02b";
			      when 174 => read_data_o <= x"d02b";
			      when 175 => read_data_o <= x"d02b";
			      when 176 => read_data_o <= x"d02b";
			      when 177 => read_data_o <= x"d02b";
			      when 178 => read_data_o <= x"d02b";
			      when 179 => read_data_o <= x"d02b";
			      when 180 => read_data_o <= x"d02b";
			      when 181 => read_data_o <= x"72c0";
			      when 182 => read_data_o <= x"0150";
			      when 183 => read_data_o <= x"d02b";
			      when 184 => read_data_o <= x"d02b";
			      when 185 => read_data_o <= x"d02b";
			      when 186 => read_data_o <= x"d02b";
			      when 187 => read_data_o <= x"d02b";
			      when 188 => read_data_o <= x"d02b";
			      when 189 => read_data_o <= x"d02b";
			      when 190 => read_data_o <= x"d02b";
			      when 191 => read_data_o <= x"72c0";
			      when 192 => read_data_o <= x"0104";
			      when 193 => read_data_o <= x"d02b";
			      when 194 => read_data_o <= x"d02b";
			      when 195 => read_data_o <= x"d02b";
			      when 196 => read_data_o <= x"d02b";
			      when 197 => read_data_o <= x"d02b";
			      when 198 => read_data_o <= x"d02b";
			      when 199 => read_data_o <= x"d02b";
			      when 200 => read_data_o <= x"d02b";
			      when 201 => read_data_o <= x"72c0";
			      when 202 => read_data_o <= x"00ec";
			      when 203 => read_data_o <= x"d02b";
			      when 204 => read_data_o <= x"d02b";
			      when 205 => read_data_o <= x"d02b";
			      when 206 => read_data_o <= x"d02b";
			      when 207 => read_data_o <= x"d02b";
			      when 208 => read_data_o <= x"d02b";
			      when 209 => read_data_o <= x"d02b";
			      when 210 => read_data_o <= x"d02b";
			      when 211 => read_data_o <= x"72c0";
			      when 212 => read_data_o <= x"00a0";
			      when 213 => read_data_o <= x"d02b";
			      when 214 => read_data_o <= x"d02b";
			      when 215 => read_data_o <= x"d02b";
			      when 216 => read_data_o <= x"d02b";
			      when 217 => read_data_o <= x"d02b";
			      when 218 => read_data_o <= x"d02b";
			      when 219 => read_data_o <= x"d02b";
			      when 220 => read_data_o <= x"d02b";
			      when 221 => read_data_o <= x"72c0";
			      when 222 => read_data_o <= x"0088";
			      when 223 => read_data_o <= x"d02b";
			      when 224 => read_data_o <= x"d02b";
			      when 225 => read_data_o <= x"d02b";
			      when 226 => read_data_o <= x"d02b";
			      when 227 => read_data_o <= x"d02b";
			      when 228 => read_data_o <= x"d02b";
			      when 229 => read_data_o <= x"d02b";
			      when 230 => read_data_o <= x"d02b";
			      when 231 => read_data_o <= x"a1d0";
			      when 232 => read_data_o <= x"72c0";
			      when 233 => read_data_o <= x"0030";
			      when 234 => read_data_o <= x"d0a1";
			      when 235 => read_data_o <= x"d095";
			      when 236 => read_data_o <= x"d1a8";
			      when 237 => read_data_o <= x"d17f";
			      when 238 => read_data_o <= x"d30c";
			      when 239 => read_data_o <= x"d1da";
			      when 240 => read_data_o <= x"d160";
			      when 241 => read_data_o <= x"d16b";
			      when 242 => read_data_o <= x"72c0";
			      when 243 => read_data_o <= x"0050";
			      when 244 => read_data_o <= x"d160";
			      when 245 => read_data_o <= x"d1da";
			      when 246 => read_data_o <= x"d1da";
			      when 247 => read_data_o <= x"d02b";
			      when 248 => read_data_o <= x"d0b2";
			      when 249 => read_data_o <= x"d0b2";
			      when 250 => read_data_o <= x"d0d1";
			      when 251 => read_data_o <= x"d02b";
			      when 252 => read_data_o <= x"2403";
			      when 253 => read_data_o <= x"7060";
			      when 254 => read_data_o <= x"01e8";
			      when 255 => read_data_o <= x"d02b";
			      when 256 => read_data_o <= x"d02b";
			      when 257 => read_data_o <= x"d02b";
			      when 258 => read_data_o <= x"d02b";
			      when 259 => read_data_o <= x"d02b";
			      when 260 => read_data_o <= x"d02b";
			      when 261 => read_data_o <= x"d02b";
			      when 262 => read_data_o <= x"d02b";
			      when 263 => read_data_o <= x"d02b";
			      when 264 => read_data_o <= x"d02b";
			      when 265 => read_data_o <= x"d02b";
			      when 266 => read_data_o <= x"d02b";
			      when 267 => read_data_o <= x"d02b";
			      when 268 => read_data_o <= x"d02b";
			      when 269 => read_data_o <= x"d02b";
			      when 270 => read_data_o <= x"d02b";
			      when 271 => read_data_o <= x"d02b";
			      when 272 => read_data_o <= x"d02b";
			      when 273 => read_data_o <= x"d02b";
			      when 274 => read_data_o <= x"d02b";
			      when 275 => read_data_o <= x"d02b";
			      when 276 => read_data_o <= x"d02b";
			      when 277 => read_data_o <= x"d02b";
			      when 278 => read_data_o <= x"d02b";
			      when 279 => read_data_o <= x"d02b";
			      when 280 => read_data_o <= x"d02b";
			      when 281 => read_data_o <= x"d02b";
			      when 282 => read_data_o <= x"d02b";
			      when 283 => read_data_o <= x"d02b";
			      when 284 => read_data_o <= x"d02b";
			      when 285 => read_data_o <= x"d02b";
			      when 286 => read_data_o <= x"d02b";
			      when 287 => read_data_o <= x"7060";
			      when 288 => read_data_o <= x"0202";
			      when 289 => read_data_o <= x"d02b";
			      when 290 => read_data_o <= x"d02b";
			      when 291 => read_data_o <= x"d02b";
			      when 292 => read_data_o <= x"d02b";
			      when 293 => read_data_o <= x"d02b";
			      when 294 => read_data_o <= x"d02b";
			      when 295 => read_data_o <= x"d02b";
			      when 296 => read_data_o <= x"d02b";
			      when 297 => read_data_o <= x"d02b";
			      when 298 => read_data_o <= x"d02b";
			      when 299 => read_data_o <= x"d02b";
			      when 300 => read_data_o <= x"d02b";
			      when 301 => read_data_o <= x"d02b";
			      when 302 => read_data_o <= x"d02b";
			      when 303 => read_data_o <= x"d02b";
			      when 304 => read_data_o <= x"d02b";
			      when 305 => read_data_o <= x"d02b";
			      when 306 => read_data_o <= x"d02b";
			      when 307 => read_data_o <= x"d02b";
			      when 308 => read_data_o <= x"d02b";
			      when 309 => read_data_o <= x"d02b";
			      when 310 => read_data_o <= x"d02b";
			      when 311 => read_data_o <= x"d02b";
			      when 312 => read_data_o <= x"d02b";
			      when 313 => read_data_o <= x"d02b";
			      when 314 => read_data_o <= x"d02b";
			      when 315 => read_data_o <= x"d02b";
			      when 316 => read_data_o <= x"d02b";
			      when 317 => read_data_o <= x"d02b";
			      when 318 => read_data_o <= x"d02b";
			      when 319 => read_data_o <= x"d02b";
			      when 320 => read_data_o <= x"d02b";
			      when 321 => read_data_o <= x"7060";
			      when 322 => read_data_o <= x"0224";
			      when 323 => read_data_o <= x"d02b";
			      when 324 => read_data_o <= x"d02b";
			      when 325 => read_data_o <= x"d02b";
			      when 326 => read_data_o <= x"d02b";
			      when 327 => read_data_o <= x"d02b";
			      when 328 => read_data_o <= x"d137";
			      when 329 => read_data_o <= x"d1a8";
			      when 330 => read_data_o <= x"d1c5";
			      when 331 => read_data_o <= x"d1a2";
			      when 332 => read_data_o <= x"d1ef";
			      when 333 => read_data_o <= x"d157";
			      when 334 => read_data_o <= x"d02b";
			      when 335 => read_data_o <= x"d157";
			      when 336 => read_data_o <= x"d137";
			      when 337 => read_data_o <= x"d1ef";
			      when 338 => read_data_o <= x"d137";
			      when 339 => read_data_o <= x"d02b";
			      when 340 => read_data_o <= x"d02b";
			      when 341 => read_data_o <= x"d02b";
			      when 342 => read_data_o <= x"7060";
			      when 343 => read_data_o <= x"023e";
			      when 344 => read_data_o <= x"d1da";
			      when 345 => read_data_o <= x"d16b";
			      when 346 => read_data_o <= x"d02b";
			      when 347 => read_data_o <= x"d137";
			      when 348 => read_data_o <= x"d157";
			      when 349 => read_data_o <= x"d191";
			      when 350 => read_data_o <= x"d1f6";
			      when 351 => read_data_o <= x"d1e5";
			      when 352 => read_data_o <= x"d1ef";
			      when 353 => read_data_o <= x"d02b";
			      when 354 => read_data_o <= x"d1e5";
			      when 355 => read_data_o <= x"d1ef";
			      when 356 => read_data_o <= x"d137";
			      when 357 => read_data_o <= x"d1ef";
			      when 358 => read_data_o <= x"d1f6";
			      when 359 => read_data_o <= x"d1e5";
			      when 360 => read_data_o <= x"d0fa";
			      when 361 => read_data_o <= x"d02b";
			      when 362 => read_data_o <= x"d02b";
			      when 363 => read_data_o <= x"71b2";
			      when 364 => read_data_o <= x"02ba";
			      when 365 => read_data_o <= x"d02b";
			      when 366 => read_data_o <= x"d02b";
			      when 367 => read_data_o <= x"d02b";
			      when 368 => read_data_o <= x"d02b";
			      when 369 => read_data_o <= x"d02b";
			      when 370 => read_data_o <= x"d02b";
			      when 371 => read_data_o <= x"d02b";
			      when 372 => read_data_o <= x"d02b";
			      when 373 => read_data_o <= x"d02b";
			      when 374 => read_data_o <= x"d02b";
			      when 375 => read_data_o <= x"d02b";
			      when 376 => read_data_o <= x"d02b";
			      when 377 => read_data_o <= x"d02b";
			      when 378 => read_data_o <= x"d02b";
			      when 379 => read_data_o <= x"d02b";
			      when 380 => read_data_o <= x"d02b";
			      when 381 => read_data_o <= x"71b2";
			      when 382 => read_data_o <= x"029c";
			      when 383 => read_data_o <= x"d02b";
			      when 384 => read_data_o <= x"d02b";
			      when 385 => read_data_o <= x"d02b";
			      when 386 => read_data_o <= x"d02b";
			      when 387 => read_data_o <= x"d02b";
			      when 388 => read_data_o <= x"d02b";
			      when 389 => read_data_o <= x"d02b";
			      when 390 => read_data_o <= x"d02b";
			      when 391 => read_data_o <= x"d02b";
			      when 392 => read_data_o <= x"d02b";
			      when 393 => read_data_o <= x"d02b";
			      when 394 => read_data_o <= x"d02b";
			      when 395 => read_data_o <= x"d02b";
			      when 396 => read_data_o <= x"d02b";
			      when 397 => read_data_o <= x"d02b";
			      when 398 => read_data_o <= x"d02b";
			      when 399 => read_data_o <= x"7040";
			      when 400 => read_data_o <= x"0030";
			      when 401 => read_data_o <= x"d02b";
			      when 402 => read_data_o <= x"d1da";
			      when 403 => read_data_o <= x"d140";
			      when 404 => read_data_o <= x"d204";
			      when 405 => read_data_o <= x"d02b";
			      when 406 => read_data_o <= x"d0a1";
			      when 407 => read_data_o <= x"d08c";
			      when 408 => read_data_o <= x"d095";
			      when 409 => read_data_o <= x"d1a8";
			      when 410 => read_data_o <= x"d17f";
			      when 411 => read_data_o <= x"d30c";
			      when 412 => read_data_o <= x"7110";
			      when 413 => read_data_o <= x"0030";
			      when 414 => read_data_o <= x"d02b";
			      when 415 => read_data_o <= x"d1fe";
			      when 416 => read_data_o <= x"d140";
			      when 417 => read_data_o <= x"d204";
			      when 418 => read_data_o <= x"d02b";
			      when 419 => read_data_o <= x"d0a1";
			      when 420 => read_data_o <= x"d08c";
			      when 421 => read_data_o <= x"d095";
			      when 422 => read_data_o <= x"d1a8";
			      when 423 => read_data_o <= x"d17f";
			      when 424 => read_data_o <= x"d30c";
			      when 425 => read_data_o <= x"71f0";
			      when 426 => read_data_o <= x"0030";
			      when 427 => read_data_o <= x"d02b";
			      when 428 => read_data_o <= x"d1e5";
			      when 429 => read_data_o <= x"d204";
			      when 430 => read_data_o <= x"d1c5";
			      when 431 => read_data_o <= x"d02b";
			      when 432 => read_data_o <= x"d0c6";
			      when 433 => read_data_o <= x"d0b2";
			      when 434 => read_data_o <= x"d095";
			      when 435 => read_data_o <= x"d2a8";
			      when 436 => read_data_o <= x"d2dc";
			      when 437 => read_data_o <= x"d02b";
			      when 438 => read_data_o <= x"d02b";
			      when 439 => read_data_o <= x"71e0";
			      when 440 => read_data_o <= x"0050";
			      when 441 => read_data_o <= x"d1e5";
			      when 442 => read_data_o <= x"d1c5";
			      when 443 => read_data_o <= x"d137";
			      when 444 => read_data_o <= x"d1b2";
			      when 445 => read_data_o <= x"d02b";
			      when 446 => read_data_o <= x"d0a8";
			      when 447 => read_data_o <= x"d0d1";
			      when 448 => read_data_o <= x"d08c";
			      when 449 => read_data_o <= x"d0c6";
			      when 450 => read_data_o <= x"d095";
			      when 451 => read_data_o <= x"d174";
			      when 452 => read_data_o <= x"d17f";
			      when 453 => read_data_o <= x"d30c";
			      when 454 => read_data_o <= x"d02b";
			      when 455 => read_data_o <= x"d02b";
			      when 456 => read_data_o <= x"d02b";
			      when 457 => read_data_o <= x"d02b";
			      when 458 => read_data_o <= x"d02b";
			      when 459 => read_data_o <= x"7050";
			      when 460 => read_data_o <= x"0050";
			      when 461 => read_data_o <= x"d14e";
			      when 462 => read_data_o <= x"d160";
			      when 463 => read_data_o <= x"d1b2";
			      when 464 => read_data_o <= x"d1ef";
			      when 465 => read_data_o <= x"d160";
			      when 466 => read_data_o <= x"d1da";
			      when 467 => read_data_o <= x"d02b";
			      when 468 => read_data_o <= x"d0a1";
			      when 469 => read_data_o <= x"d0b2";
			      when 470 => read_data_o <= x"d08c";
			      when 471 => read_data_o <= x"d0a8";
			      when 472 => read_data_o <= x"d0c6";
			      when 473 => read_data_o <= x"d174";
			      when 474 => read_data_o <= x"d17f";
			      when 475 => read_data_o <= x"d30c";
			      when 476 => read_data_o <= x"d02b";
			      when 477 => read_data_o <= x"d02b";
			      when 478 => read_data_o <= x"d02b";
			      when 479 => read_data_o <= x"d02b";
			      when 480 => read_data_o <= x"d02b";
			      when 481 => read_data_o <= x"d02b";
			      when 482 => read_data_o <= x"d02b";
			      when 483 => read_data_o <= x"7050";
			      when 484 => read_data_o <= x"02dc";
			      when 485 => read_data_o <= x"d1da";
			      when 486 => read_data_o <= x"d1a2";
			      when 487 => read_data_o <= x"d02b";
			      when 488 => read_data_o <= x"d095";
			      when 489 => read_data_o <= x"d25f";
			      when 490 => read_data_o <= x"d140";
			      when 491 => read_data_o <= x"d2a8";
			      when 492 => read_data_o <= x"d02b";
			      when 493 => read_data_o <= x"d02b";
			      when 494 => read_data_o <= x"d02b";
			      when 495 => read_data_o <= x"d02b";
			      when 496 => read_data_o <= x"d02b";
			      when 497 => read_data_o <= x"d02b";
			      when 498 => read_data_o <= x"7040";
			      when 499 => read_data_o <= x"02fc";
			      when 500 => read_data_o <= x"d02b";
			      when 501 => read_data_o <= x"d137";
			      when 502 => read_data_o <= x"d1ef";
			      when 503 => read_data_o <= x"d1ef";
			      when 504 => read_data_o <= x"d160";
			      when 505 => read_data_o <= x"d1b2";
			      when 506 => read_data_o <= x"d02b";
			      when 507 => read_data_o <= x"d0a1";
			      when 508 => read_data_o <= x"d095";
			      when 509 => read_data_o <= x"d25f";
			      when 510 => read_data_o <= x"d140";
			      when 511 => read_data_o <= x"7110";
			      when 512 => read_data_o <= x"02fc";
			      when 513 => read_data_o <= x"d02b";
			      when 514 => read_data_o <= x"d02b";
			      when 515 => read_data_o <= x"d02b";
			      when 516 => read_data_o <= x"d02b";
			      when 517 => read_data_o <= x"d02b";
			      when 518 => read_data_o <= x"d02b";
			      when 519 => read_data_o <= x"d02b";
			      when 520 => read_data_o <= x"d02b";
			      when 521 => read_data_o <= x"7130";
			      when 522 => read_data_o <= x"02dc";
			      when 523 => read_data_o <= x"d0a1";
			      when 524 => read_data_o <= x"d095";
			      when 525 => read_data_o <= x"d25f";
			      when 526 => read_data_o <= x"d140";
			      when 527 => read_data_o <= x"d091";
			      when 528 => read_data_o <= x"d02b";
			      when 529 => read_data_o <= x"71b0";
			      when 530 => read_data_o <= x"02fc";
			      when 531 => read_data_o <= x"d02b";
			      when 532 => read_data_o <= x"d02b";
			      when 533 => read_data_o <= x"d02b";
			      when 534 => read_data_o <= x"d02b";
			      when 535 => read_data_o <= x"d02b";
			      when 536 => read_data_o <= x"d02b";
			      when 537 => read_data_o <= x"d02b";
			      when 538 => read_data_o <= x"d02b";
			      when 539 => read_data_o <= x"d02b";
			      when 540 => read_data_o <= x"d02b";
			      when 541 => read_data_o <= x"d02b";
			      when 542 => read_data_o <= x"d02b";
			      when 543 => read_data_o <= x"d02b";
			      when 544 => read_data_o <= x"d02b";
			      when 545 => read_data_o <= x"d02b";
			      when 546 => read_data_o <= x"d02b";
			      when 547 => read_data_o <= x"d02b";
			      when 548 => read_data_o <= x"71b0";
			      when 549 => read_data_o <= x"02dc";
			      when 550 => read_data_o <= x"d02b";
			      when 551 => read_data_o <= x"d02b";
			      when 552 => read_data_o <= x"d02b";
			      when 553 => read_data_o <= x"d02b";
			      when 554 => read_data_o <= x"d02b";
			      when 555 => read_data_o <= x"d02b";
			      when 556 => read_data_o <= x"d02b";
			      when 557 => read_data_o <= x"d02b";
			      when 558 => read_data_o <= x"d02b";
			      when 559 => read_data_o <= x"d02b";
			      when 560 => read_data_o <= x"d02b";
			      when 561 => read_data_o <= x"d02b";
			      when 562 => read_data_o <= x"d02b";
			      when 563 => read_data_o <= x"d02b";
			      when 564 => read_data_o <= x"d02b";
			      when 565 => read_data_o <= x"d02b";
			      when 566 => read_data_o <= x"d02b";
			      when 567 => read_data_o <= x"d02b";
			      when 568 => read_data_o <= x"d02b";
			      when 569 => read_data_o <= x"7060";
			      when 570 => read_data_o <= x"027a";
			      when 571 => read_data_o <= x"d02b";
			      when 572 => read_data_o <= x"d02b";
			      when 573 => read_data_o <= x"d02b";
			      when 574 => read_data_o <= x"d02b";
			      when 575 => read_data_o <= x"d02b";
			      when 576 => read_data_o <= x"d02b";
			      when 577 => read_data_o <= x"d02b";
			      when 578 => read_data_o <= x"d02b";
			      when 579 => read_data_o <= x"d02b";
			      when 580 => read_data_o <= x"d02b";
			      when 581 => read_data_o <= x"d02b";
			      when 582 => read_data_o <= x"d02b";
			      when 583 => read_data_o <= x"7040";
			      when 584 => read_data_o <= x"022c";
			      when 585 => read_data_o <= x"d02b";
			      when 586 => read_data_o <= x"7040";
			      when 587 => read_data_o <= x"020c";
			      when 588 => read_data_o <= x"d02b";
			      when 589 => read_data_o <= x"7040";
			      when 590 => read_data_o <= x"01ec";
			      when 591 => read_data_o <= x"d02b";
			      when 592 => read_data_o <= x"7040";
			      when 593 => read_data_o <= x"01cc";
			      when 594 => read_data_o <= x"d02b";
			      when 595 => read_data_o <= x"7040";
			      when 596 => read_data_o <= x"01ac";
			      when 597 => read_data_o <= x"d02b";
			      when 598 => read_data_o <= x"7040";
			      when 599 => read_data_o <= x"018c";
			      when 600 => read_data_o <= x"d02b";
			      when 601 => read_data_o <= x"7040";
			      when 602 => read_data_o <= x"016c";
			      when 603 => read_data_o <= x"d02b";
			      when 604 => read_data_o <= x"7040";
			      when 605 => read_data_o <= x"014c";
			      when 606 => read_data_o <= x"d02b";
			      when 607 => read_data_o <= x"7040";
			      when 608 => read_data_o <= x"012c";
			      when 609 => read_data_o <= x"d02b";
			      when 610 => read_data_o <= x"7040";
			      when 611 => read_data_o <= x"010c";
			      when 612 => read_data_o <= x"d02b";
			      when 613 => read_data_o <= x"ba04";
			      when 614 => read_data_o <= x"a000";
			      when 615 => read_data_o <= x"a000";
			      when 616 => read_data_o <= x"7290";
			      when 617 => read_data_o <= x"0270";
			      when 618 => read_data_o <= x"d074";
			      when 619 => read_data_o <= x"2404";
			      when 620 => read_data_o <= x"7064";
			      when 621 => read_data_o <= x"02bc";
			      when 622 => read_data_o <= x"a532";
			      when 623 => read_data_o <= x"a000";
			      when 624 => read_data_o <= x"a000";
			      when 625 => read_data_o <= x"a000";
			      when 626 => read_data_o <= x"a000";
			      when 627 => read_data_o <= x"a000";
			      when 628 => read_data_o <= x"a000";
			      when 629 => read_data_o <= x"a000";
			      when 630 => read_data_o <= x"a000";
			      when 631 => read_data_o <= x"a000";
			      when 632 => read_data_o <= x"a000";
			      when 633 => read_data_o <= x"a000";
			      when 634 => read_data_o <= x"a000";
			      when 635 => read_data_o <= x"a000";
			      when 636 => read_data_o <= x"a000";
			      when 637 => read_data_o <= x"a000";
			      when 638 => read_data_o <= x"a000";
			      when 639 => read_data_o <= x"a000";
			      when 640 => read_data_o <= x"a000";
			      when 641 => read_data_o <= x"a000";
			      when 642 => read_data_o <= x"a000";
			      when 643 => read_data_o <= x"a000";
			      when 644 => read_data_o <= x"a000";
			      when 645 => read_data_o <= x"a000";
			      when 646 => read_data_o <= x"a000";
			      when 647 => read_data_o <= x"a000";
			      when 648 => read_data_o <= x"a000";
			      when 649 => read_data_o <= x"a000";
			      when 650 => read_data_o <= x"a000";
			      when 651 => read_data_o <= x"a000";
			      when 652 => read_data_o <= x"a000";
			      when 653 => read_data_o <= x"a000";
			      when 654 => read_data_o <= x"a000";
			      when 655 => read_data_o <= x"a000";
			      when 656 => read_data_o <= x"a000";
			      when 657 => read_data_o <= x"a000";
			      when 658 => read_data_o <= x"a000";
			      when 659 => read_data_o <= x"a000";
			      when 660 => read_data_o <= x"a000";
			      when 661 => read_data_o <= x"a000";
			      when 662 => read_data_o <= x"a000";
			      when 663 => read_data_o <= x"a000";
			      when 664 => read_data_o <= x"a000";
			      when 665 => read_data_o <= x"2403";
			      when 666 => read_data_o <= x"7064";
			      when 667 => read_data_o <= x"02bc";
when 668 => read_data_o <= x"a58e";
when 669 => read_data_o <= x"a000";
when 670 => read_data_o <= x"a000";
when 671 => read_data_o <= x"a000";
when 672 => read_data_o <= x"a000";
when 673 => read_data_o <= x"a000";
when 674 => read_data_o <= x"a000";
when 675 => read_data_o <= x"a000";
when 676 => read_data_o <= x"a000";
when 677 => read_data_o <= x"a000";
when 678 => read_data_o <= x"a000";
when 679 => read_data_o <= x"a000";
when 680 => read_data_o <= x"a000";
when 681 => read_data_o <= x"a000";
when 682 => read_data_o <= x"a000";
when 683 => read_data_o <= x"a000";
when 684 => read_data_o <= x"a000";
when 685 => read_data_o <= x"a000";
when 686 => read_data_o <= x"a000";
when 687 => read_data_o <= x"a000";
when 688 => read_data_o <= x"a000";
when 689 => read_data_o <= x"a000";
when 690 => read_data_o <= x"a000";
when 691 => read_data_o <= x"a000";
when 692 => read_data_o <= x"a000";
when 693 => read_data_o <= x"a000";
when 694 => read_data_o <= x"a000";
when 695 => read_data_o <= x"a000";
when 696 => read_data_o <= x"a000";
when 697 => read_data_o <= x"a000";
when 698 => read_data_o <= x"a000";
when 699 => read_data_o <= x"a000";
when 700 => read_data_o <= x"a000";
when 701 => read_data_o <= x"a000";
when 702 => read_data_o <= x"a000";
when 703 => read_data_o <= x"a000";
when 704 => read_data_o <= x"a000";
when 705 => read_data_o <= x"a000";
when 706 => read_data_o <= x"a000";
when 707 => read_data_o <= x"a000";
when 708 => read_data_o <= x"a000";
when 709 => read_data_o <= x"a000";
when 710 => read_data_o <= x"a000";
when 711 => read_data_o <= x"2401";
when 712 => read_data_o <= x"a592";
when 713 => read_data_o <= x"7064";
when 714 => read_data_o <= x"0064";
when 715 => read_data_o <= x"7064";
when 716 => read_data_o <= x"0064";
when 717 => read_data_o <= x"5064";
when 718 => read_data_o <= x"0190";
when 719 => read_data_o <= x"5064";
when 720 => read_data_o <= x"02bc";
when 721 => read_data_o <= x"70a0";
when 722 => read_data_o <= x"02bc";
when 723 => read_data_o <= x"50a0";
when 724 => read_data_o <= x"0190";
when 725 => read_data_o <= x"50a0";
when 726 => read_data_o <= x"0064";
when 727 => read_data_o <= x"70dc";
when 728 => read_data_o <= x"0064";
when 729 => read_data_o <= x"50dc";
when 730 => read_data_o <= x"0190";
when 731 => read_data_o <= x"50dc";
when 732 => read_data_o <= x"02bc";
when 733 => read_data_o <= x"7118";
when 734 => read_data_o <= x"02bc";
when 735 => read_data_o <= x"5118";
when 736 => read_data_o <= x"0190";
when 737 => read_data_o <= x"5118";
when 738 => read_data_o <= x"0064";
when 739 => read_data_o <= x"7154";
when 740 => read_data_o <= x"0064";
when 741 => read_data_o <= x"5154";
when 742 => read_data_o <= x"0190";
when 743 => read_data_o <= x"5154";
when 744 => read_data_o <= x"02bc";
when 745 => read_data_o <= x"7190";
when 746 => read_data_o <= x"02bc";
when 747 => read_data_o <= x"5190";
when 748 => read_data_o <= x"0190";
when 749 => read_data_o <= x"5190";
when 750 => read_data_o <= x"0064";
when 751 => read_data_o <= x"71cc";
when 752 => read_data_o <= x"0064";
when 753 => read_data_o <= x"51cc";
when 754 => read_data_o <= x"0190";
when 755 => read_data_o <= x"51cc";
when 756 => read_data_o <= x"02bc";
when 757 => read_data_o <= x"7208";
when 758 => read_data_o <= x"02bc";
when 759 => read_data_o <= x"5208";
when 760 => read_data_o <= x"0190";
when 761 => read_data_o <= x"5208";
when 762 => read_data_o <= x"0064";
when 763 => read_data_o <= x"7244";
when 764 => read_data_o <= x"0064";
when 765 => read_data_o <= x"5244";
when 766 => read_data_o <= x"0190";
when 767 => read_data_o <= x"5244";
when 768 => read_data_o <= x"02bc";
when 769 => read_data_o <= x"7280";
when 770 => read_data_o <= x"02bc";
when 771 => read_data_o <= x"5280";
when 772 => read_data_o <= x"0190";
when 773 => read_data_o <= x"5280";
when 774 => read_data_o <= x"0064";
when 775 => read_data_o <= x"72bc";
when 776 => read_data_o <= x"0064";
when 777 => read_data_o <= x"52bc";
when 778 => read_data_o <= x"0190";
when 779 => read_data_o <= x"52bc";
when 780 => read_data_o <= x"02bc";
when 781 => read_data_o <= x"72bc";
when 782 => read_data_o <= x"02bc";
when 783 => read_data_o <= x"5190";
when 784 => read_data_o <= x"02bc";
when 785 => read_data_o <= x"5064";
when 786 => read_data_o <= x"02bc";
when 787 => read_data_o <= x"7064";
when 788 => read_data_o <= x"0280";
when 789 => read_data_o <= x"5190";
when 790 => read_data_o <= x"0280";
when 791 => read_data_o <= x"52bc";
when 792 => read_data_o <= x"0280";
when 793 => read_data_o <= x"72bc";
when 794 => read_data_o <= x"0244";
when 795 => read_data_o <= x"5190";
when 796 => read_data_o <= x"0244";
when 797 => read_data_o <= x"5064";
when 798 => read_data_o <= x"0244";
when 799 => read_data_o <= x"7064";
when 800 => read_data_o <= x"0208";
when 801 => read_data_o <= x"5190";
when 802 => read_data_o <= x"0208";
when 803 => read_data_o <= x"52bc";
when 804 => read_data_o <= x"0208";
when 805 => read_data_o <= x"72bc";
when 806 => read_data_o <= x"01cc";
when 807 => read_data_o <= x"5190";
when 808 => read_data_o <= x"01cc";
when 809 => read_data_o <= x"5064";
when 810 => read_data_o <= x"01cc";
when 811 => read_data_o <= x"7064";
when 812 => read_data_o <= x"0190";
when 813 => read_data_o <= x"5190";
when 814 => read_data_o <= x"0190";
when 815 => read_data_o <= x"52bc";
when 816 => read_data_o <= x"0190";
when 817 => read_data_o <= x"72bc";
when 818 => read_data_o <= x"0154";
when 819 => read_data_o <= x"5190";
when 820 => read_data_o <= x"0154";
when 821 => read_data_o <= x"5064";
when 822 => read_data_o <= x"0154";
when 823 => read_data_o <= x"7064";
when 824 => read_data_o <= x"0118";
when 825 => read_data_o <= x"5190";
when 826 => read_data_o <= x"0118";
when 827 => read_data_o <= x"52bc";
when 828 => read_data_o <= x"0118";
when 829 => read_data_o <= x"72bc";
when 830 => read_data_o <= x"00dc";
when 831 => read_data_o <= x"5190";
when 832 => read_data_o <= x"00dc";
when 833 => read_data_o <= x"5064";
when 834 => read_data_o <= x"00dc";
when 835 => read_data_o <= x"7064";
when 836 => read_data_o <= x"00a0";
when 837 => read_data_o <= x"5190";
when 838 => read_data_o <= x"00a0";
when 839 => read_data_o <= x"52bc";
when 840 => read_data_o <= x"00a0";
when 841 => read_data_o <= x"72bc";
when 842 => read_data_o <= x"0064";
when 843 => read_data_o <= x"5190";
when 844 => read_data_o <= x"0064";
when 845 => read_data_o <= x"5064";
when 846 => read_data_o <= x"0064";
when 847 => read_data_o <= x"a6a0";
when 848 => read_data_o <= x"2403";
when 849 => read_data_o <= x"a6e2";
when 850 => read_data_o <= x"a000";
when 851 => read_data_o <= x"a000";
when 852 => read_data_o <= x"a000";
when 853 => read_data_o <= x"a000";
when 854 => read_data_o <= x"a000";
when 855 => read_data_o <= x"a000";
when 856 => read_data_o <= x"a000";
when 857 => read_data_o <= x"a000";
when 858 => read_data_o <= x"a000";
when 859 => read_data_o <= x"a000";
when 860 => read_data_o <= x"a000";
when 861 => read_data_o <= x"a000";
when 862 => read_data_o <= x"a000";
when 863 => read_data_o <= x"a000";
when 864 => read_data_o <= x"a000";
when 865 => read_data_o <= x"a000";
when 866 => read_data_o <= x"a000";
when 867 => read_data_o <= x"a000";
when 868 => read_data_o <= x"a000";
when 869 => read_data_o <= x"a000";
when 870 => read_data_o <= x"a000";
when 871 => read_data_o <= x"a000";
when 872 => read_data_o <= x"a000";
when 873 => read_data_o <= x"a000";
when 874 => read_data_o <= x"a000";
when 875 => read_data_o <= x"a000";
when 876 => read_data_o <= x"a000";
when 877 => read_data_o <= x"a000";
when 878 => read_data_o <= x"a000";
when 879 => read_data_o <= x"a000";
when 880 => read_data_o <= x"a000";
when 881 => read_data_o <= x"a722";
when 882 => read_data_o <= x"a000";
when 883 => read_data_o <= x"a000";
when 884 => read_data_o <= x"a000";
when 885 => read_data_o <= x"a000";
when 886 => read_data_o <= x"a000";
when 887 => read_data_o <= x"a000";
when 888 => read_data_o <= x"a000";
when 889 => read_data_o <= x"a000";
when 890 => read_data_o <= x"a000";
when 891 => read_data_o <= x"a000";
when 892 => read_data_o <= x"a000";
when 893 => read_data_o <= x"a000";
when 894 => read_data_o <= x"a000";
when 895 => read_data_o <= x"a000";
when 896 => read_data_o <= x"a000";
when 897 => read_data_o <= x"a000";
when 898 => read_data_o <= x"a000";
when 899 => read_data_o <= x"a000";
when 900 => read_data_o <= x"a000";
when 901 => read_data_o <= x"a000";
when 902 => read_data_o <= x"a000";
when 903 => read_data_o <= x"a000";
when 904 => read_data_o <= x"a000";
when 905 => read_data_o <= x"a000";
when 906 => read_data_o <= x"a000";
when 907 => read_data_o <= x"a000";
when 908 => read_data_o <= x"a000";
when 909 => read_data_o <= x"a000";
when 910 => read_data_o <= x"a000";
when 911 => read_data_o <= x"a000";
when 912 => read_data_o <= x"a000";
when 913 => read_data_o <= x"a762";
when 914 => read_data_o <= x"a000";
when 915 => read_data_o <= x"a000";
when 916 => read_data_o <= x"a000";
when 917 => read_data_o <= x"a000";
when 918 => read_data_o <= x"a000";
when 919 => read_data_o <= x"a000";
when 920 => read_data_o <= x"a000";
when 921 => read_data_o <= x"a000";
when 922 => read_data_o <= x"a000";
when 923 => read_data_o <= x"a000";
when 924 => read_data_o <= x"a000";
when 925 => read_data_o <= x"a000";
when 926 => read_data_o <= x"a000";
when 927 => read_data_o <= x"a000";
when 928 => read_data_o <= x"a000";
when 929 => read_data_o <= x"a000";
when 930 => read_data_o <= x"a000";
when 931 => read_data_o <= x"a000";
when 932 => read_data_o <= x"a000";
when 933 => read_data_o <= x"a000";
when 934 => read_data_o <= x"a000";
when 935 => read_data_o <= x"a000";
when 936 => read_data_o <= x"a000";
when 937 => read_data_o <= x"a000";
when 938 => read_data_o <= x"a000";
when 939 => read_data_o <= x"a000";
when 940 => read_data_o <= x"a000";
when 941 => read_data_o <= x"a000";
when 942 => read_data_o <= x"a000";
when 943 => read_data_o <= x"a000";
when 944 => read_data_o <= x"a000";
when 945 => read_data_o <= x"a7a2";
when 946 => read_data_o <= x"a000";
when 947 => read_data_o <= x"a000";
when 948 => read_data_o <= x"a000";
when 949 => read_data_o <= x"a000";
when 950 => read_data_o <= x"a000";
when 951 => read_data_o <= x"a000";
when 952 => read_data_o <= x"a000";
when 953 => read_data_o <= x"a000";
when 954 => read_data_o <= x"a000";
when 955 => read_data_o <= x"a000";
when 956 => read_data_o <= x"a000";
when 957 => read_data_o <= x"a000";
when 958 => read_data_o <= x"a000";
when 959 => read_data_o <= x"a000";
when 960 => read_data_o <= x"a000";
when 961 => read_data_o <= x"a000";
when 962 => read_data_o <= x"a000";
when 963 => read_data_o <= x"a000";
when 964 => read_data_o <= x"a000";
when 965 => read_data_o <= x"a000";
when 966 => read_data_o <= x"a000";
when 967 => read_data_o <= x"a000";
when 968 => read_data_o <= x"a000";
when 969 => read_data_o <= x"a000";
when 970 => read_data_o <= x"a000";
when 971 => read_data_o <= x"a000";
when 972 => read_data_o <= x"a000";
when 973 => read_data_o <= x"a000";
when 974 => read_data_o <= x"a000";
when 975 => read_data_o <= x"a000";
when 976 => read_data_o <= x"a000";
when 977 => read_data_o <= x"a7e2";
when 978 => read_data_o <= x"a000";
when 979 => read_data_o <= x"a000";
when 980 => read_data_o <= x"a000";
when 981 => read_data_o <= x"a000";
when 982 => read_data_o <= x"a000";
when 983 => read_data_o <= x"a000";
when 984 => read_data_o <= x"a000";
when 985 => read_data_o <= x"a000";
when 986 => read_data_o <= x"a000";
when 987 => read_data_o <= x"a000";
when 988 => read_data_o <= x"a000";
when 989 => read_data_o <= x"a000";
when 990 => read_data_o <= x"a000";
when 991 => read_data_o <= x"a000";
when 992 => read_data_o <= x"a000";
when 993 => read_data_o <= x"a000";
when 994 => read_data_o <= x"a000";
when 995 => read_data_o <= x"a000";
when 996 => read_data_o <= x"a000";
when 997 => read_data_o <= x"a000";
when 998 => read_data_o <= x"a000";
when 999 => read_data_o <= x"a000";
when 1000 => read_data_o <= x"a000";
when 1001 => read_data_o <= x"a000";
when 1002 => read_data_o <= x"a000";
when 1003 => read_data_o <= x"a000";
when 1004 => read_data_o <= x"a000";
when 1005 => read_data_o <= x"a000";
when 1006 => read_data_o <= x"a000";
when 1007 => read_data_o <= x"a000";
when 1008 => read_data_o <= x"a000";
when 1009 => read_data_o <= x"2402";
when 1010 => read_data_o <= x"7064";
when 1011 => read_data_o <= x"0064";
when 1012 => read_data_o <= x"0064";
when 1013 => read_data_o <= x"0064";
when 1014 => read_data_o <= x"0064";
when 1015 => read_data_o <= x"0064";
when 1016 => read_data_o <= x"0064";
when 1017 => read_data_o <= x"0064";
when 1018 => read_data_o <= x"0064";
when 1019 => read_data_o <= x"0064";
when 1020 => read_data_o <= x"0064";
when 1021 => read_data_o <= x"0064";
when 1022 => read_data_o <= x"0064";
when 1023 => read_data_o <= x"0064";
when 1024 => read_data_o <= x"0064";
when 1025 => read_data_o <= x"0064";
when 1026 => read_data_o <= x"0064";
when 1027 => read_data_o <= x"0064";
when 1028 => read_data_o <= x"0064";
when 1029 => read_data_o <= x"0064";
when 1030 => read_data_o <= x"0064";
when 1031 => read_data_o <= x"0064";
when 1032 => read_data_o <= x"0064";
when 1033 => read_data_o <= x"0064";
when 1034 => read_data_o <= x"0064";
when 1035 => read_data_o <= x"0064";
when 1036 => read_data_o <= x"0064";
when 1037 => read_data_o <= x"0064";
when 1038 => read_data_o <= x"0064";
when 1039 => read_data_o <= x"0064";
when 1040 => read_data_o <= x"0064";
when 1041 => read_data_o <= x"0064";
when 1042 => read_data_o <= x"0064";
when 1043 => read_data_o <= x"0064";
when 1044 => read_data_o <= x"0064";
when 1045 => read_data_o <= x"0064";
when 1046 => read_data_o <= x"0064";
when 1047 => read_data_o <= x"0064";
when 1048 => read_data_o <= x"0064";
when 1049 => read_data_o <= x"0064";
when 1050 => read_data_o <= x"0064";
when 1051 => read_data_o <= x"0064";
when 1052 => read_data_o <= x"0064";
when 1053 => read_data_o <= x"0064";
when 1054 => read_data_o <= x"0064";
when 1055 => read_data_o <= x"0064";
when 1056 => read_data_o <= x"0064";
when 1057 => read_data_o <= x"0064";
when 1058 => read_data_o <= x"0064";
when 1059 => read_data_o <= x"0064";
when 1060 => read_data_o <= x"0064";
when 1061 => read_data_o <= x"0064";
when 1062 => read_data_o <= x"0064";
when 1063 => read_data_o <= x"0064";
when 1064 => read_data_o <= x"0064";
when 1065 => read_data_o <= x"0064";
when 1066 => read_data_o <= x"0064";
when 1067 => read_data_o <= x"0064";
when 1068 => read_data_o <= x"0064";
when 1069 => read_data_o <= x"0064";
when 1070 => read_data_o <= x"0064";
when 1071 => read_data_o <= x"0064";
when 1072 => read_data_o <= x"0064";
when 1073 => read_data_o <= x"0064";
when 1074 => read_data_o <= x"0064";
when 1075 => read_data_o <= x"0064";
when 1076 => read_data_o <= x"0064";
when 1077 => read_data_o <= x"0064";
when 1078 => read_data_o <= x"0064";
when 1079 => read_data_o <= x"0064";
when 1080 => read_data_o <= x"0064";
when 1081 => read_data_o <= x"0064";
when 1082 => read_data_o <= x"0064";
when 1083 => read_data_o <= x"0064";
when 1084 => read_data_o <= x"0064";
when 1085 => read_data_o <= x"0064";
when 1086 => read_data_o <= x"0064";
when 1087 => read_data_o <= x"0064";
when 1088 => read_data_o <= x"0064";
when 1089 => read_data_o <= x"0064";
when 1090 => read_data_o <= x"0064";
when 1091 => read_data_o <= x"0064";
when 1092 => read_data_o <= x"0064";
when 1093 => read_data_o <= x"0064";
when 1094 => read_data_o <= x"0064";
when 1095 => read_data_o <= x"0064";
when 1096 => read_data_o <= x"0064";
when 1097 => read_data_o <= x"0064";
when 1098 => read_data_o <= x"0064";
when 1099 => read_data_o <= x"0064";
when 1100 => read_data_o <= x"0064";
when 1101 => read_data_o <= x"0064";
when 1102 => read_data_o <= x"0064";
when 1103 => read_data_o <= x"0064";
when 1104 => read_data_o <= x"0064";
when 1105 => read_data_o <= x"0064";
when 1106 => read_data_o <= x"0064";
when 1107 => read_data_o <= x"0064";
when 1108 => read_data_o <= x"0064";
when 1109 => read_data_o <= x"0064";
when 1110 => read_data_o <= x"0064";
when 1111 => read_data_o <= x"0064";
when 1112 => read_data_o <= x"0064";
when 1113 => read_data_o <= x"0064";
when 1114 => read_data_o <= x"0064";
when 1115 => read_data_o <= x"0064";
when 1116 => read_data_o <= x"0064";
when 1117 => read_data_o <= x"0064";
when 1118 => read_data_o <= x"0064";
when 1119 => read_data_o <= x"0064";
when 1120 => read_data_o <= x"0064";
when 1121 => read_data_o <= x"0064";
when 1122 => read_data_o <= x"0064";
when 1123 => read_data_o <= x"0064";
when 1124 => read_data_o <= x"0064";
when 1125 => read_data_o <= x"0064";
when 1126 => read_data_o <= x"0064";
when 1127 => read_data_o <= x"0064";
when 1128 => read_data_o <= x"0064";
when 1129 => read_data_o <= x"0064";
when 1130 => read_data_o <= x"0064";
when 1131 => read_data_o <= x"0064";
when 1132 => read_data_o <= x"0064";
when 1133 => read_data_o <= x"0064";
when 1134 => read_data_o <= x"0064";
when 1135 => read_data_o <= x"0064";
when 1136 => read_data_o <= x"0064";
when 1137 => read_data_o <= x"0064";
when 1138 => read_data_o <= x"0064";
when 1139 => read_data_o <= x"0064";
when 1140 => read_data_o <= x"0064";
when 1141 => read_data_o <= x"0064";
when 1142 => read_data_o <= x"0064";
when 1143 => read_data_o <= x"0064";
when 1144 => read_data_o <= x"0064";
when 1145 => read_data_o <= x"0064";
when 1146 => read_data_o <= x"0064";
when 1147 => read_data_o <= x"0064";
when 1148 => read_data_o <= x"0064";
when 1149 => read_data_o <= x"0064";
when 1150 => read_data_o <= x"0064";
when 1151 => read_data_o <= x"0064";
when 1152 => read_data_o <= x"0064";
when 1153 => read_data_o <= x"0064";
when 1154 => read_data_o <= x"0064";
when 1155 => read_data_o <= x"0064";
when 1156 => read_data_o <= x"0064";
when 1157 => read_data_o <= x"0064";
when 1158 => read_data_o <= x"0064";
when 1159 => read_data_o <= x"0064";
when 1160 => read_data_o <= x"0064";
when 1161 => read_data_o <= x"0064";
when 1162 => read_data_o <= x"0064";
when 1163 => read_data_o <= x"0064";
when 1164 => read_data_o <= x"0064";
when 1165 => read_data_o <= x"0064";
when 1166 => read_data_o <= x"0064";
when 1167 => read_data_o <= x"0064";
when 1168 => read_data_o <= x"0064";
when 1169 => read_data_o <= x"0064";
when 1170 => read_data_o <= x"0064";
when 1171 => read_data_o <= x"0064";
when 1172 => read_data_o <= x"0064";
when 1173 => read_data_o <= x"0064";
when 1174 => read_data_o <= x"0064";
when 1175 => read_data_o <= x"0064";
when 1176 => read_data_o <= x"0064";
when 1177 => read_data_o <= x"0064";
when 1178 => read_data_o <= x"0064";
when 1179 => read_data_o <= x"0064";
when 1180 => read_data_o <= x"0064";
when 1181 => read_data_o <= x"0064";
when 1182 => read_data_o <= x"0064";
when 1183 => read_data_o <= x"0064";
when 1184 => read_data_o <= x"0064";
when 1185 => read_data_o <= x"0064";
when 1186 => read_data_o <= x"0064";
when 1187 => read_data_o <= x"0064";
when 1188 => read_data_o <= x"0064";
when 1189 => read_data_o <= x"0064";
when 1190 => read_data_o <= x"0064";
when 1191 => read_data_o <= x"0064";
when 1192 => read_data_o <= x"0064";
when 1193 => read_data_o <= x"0064";
when 1194 => read_data_o <= x"0064";
when 1195 => read_data_o <= x"0064";
when 1196 => read_data_o <= x"0064";
when 1197 => read_data_o <= x"0064";
when 1198 => read_data_o <= x"0064";
when 1199 => read_data_o <= x"0064";
when 1200 => read_data_o <= x"0064";
when 1201 => read_data_o <= x"0064";
when 1202 => read_data_o <= x"0064";
when 1203 => read_data_o <= x"0064";
when 1204 => read_data_o <= x"0064";
when 1205 => read_data_o <= x"0064";
when 1206 => read_data_o <= x"0064";
when 1207 => read_data_o <= x"0064";
when 1208 => read_data_o <= x"0064";
when 1209 => read_data_o <= x"0064";
when 1210 => read_data_o <= x"0064";
when 1211 => read_data_o <= x"0064";
when 1212 => read_data_o <= x"0064";
when 1213 => read_data_o <= x"0064";
when 1214 => read_data_o <= x"0064";
when 1215 => read_data_o <= x"0064";
when 1216 => read_data_o <= x"0064";
when 1217 => read_data_o <= x"0064";
when 1218 => read_data_o <= x"0064";
when 1219 => read_data_o <= x"0064";
when 1220 => read_data_o <= x"0064";
when 1221 => read_data_o <= x"0064";
when 1222 => read_data_o <= x"0064";
when 1223 => read_data_o <= x"0064";
when 1224 => read_data_o <= x"0064";
when 1225 => read_data_o <= x"0064";
when 1226 => read_data_o <= x"0064";
when 1227 => read_data_o <= x"0064";
when 1228 => read_data_o <= x"0064";
when 1229 => read_data_o <= x"0064";
when 1230 => read_data_o <= x"0064";
when 1231 => read_data_o <= x"0064";
when 1232 => read_data_o <= x"0064";
when 1233 => read_data_o <= x"0064";
when 1234 => read_data_o <= x"0064";
when 1235 => read_data_o <= x"0064";
when 1236 => read_data_o <= x"0064";
when 1237 => read_data_o <= x"0064";
when 1238 => read_data_o <= x"0064";
when 1239 => read_data_o <= x"0064";
when 1240 => read_data_o <= x"0064";
when 1241 => read_data_o <= x"0064";
when 1242 => read_data_o <= x"0064";
when 1243 => read_data_o <= x"0064";
when 1244 => read_data_o <= x"0064";
when 1245 => read_data_o <= x"0064";
when 1246 => read_data_o <= x"0064";
when 1247 => read_data_o <= x"0064";
when 1248 => read_data_o <= x"0064";
when 1249 => read_data_o <= x"0064";
when 1250 => read_data_o <= x"0064";
when 1251 => read_data_o <= x"0064";
when 1252 => read_data_o <= x"0064";
when 1253 => read_data_o <= x"0064";
when 1254 => read_data_o <= x"0064";
when 1255 => read_data_o <= x"0064";
when 1256 => read_data_o <= x"0064";
when 1257 => read_data_o <= x"0064";
when 1258 => read_data_o <= x"0064";
when 1259 => read_data_o <= x"0064";
when 1260 => read_data_o <= x"0064";
when 1261 => read_data_o <= x"0064";
when 1262 => read_data_o <= x"0064";
when 1263 => read_data_o <= x"0064";
when 1264 => read_data_o <= x"0064";
when 1265 => read_data_o <= x"0064";
when 1266 => read_data_o <= x"0064";
when 1267 => read_data_o <= x"0064";
when 1268 => read_data_o <= x"0064";
when 1269 => read_data_o <= x"0064";
when 1270 => read_data_o <= x"0064";
when 1271 => read_data_o <= x"0064";
when 1272 => read_data_o <= x"0064";
when 1273 => read_data_o <= x"0064";
when 1274 => read_data_o <= x"0064";
when 1275 => read_data_o <= x"0064";
when 1276 => read_data_o <= x"0064";
when 1277 => read_data_o <= x"0064";
when 1278 => read_data_o <= x"0064";
when 1279 => read_data_o <= x"0064";
when 1280 => read_data_o <= x"0064";
when 1281 => read_data_o <= x"0064";
when 1282 => read_data_o <= x"0064";
when 1283 => read_data_o <= x"0064";
when 1284 => read_data_o <= x"0064";
when 1285 => read_data_o <= x"0064";
when 1286 => read_data_o <= x"0064";
when 1287 => read_data_o <= x"0064";
when 1288 => read_data_o <= x"0064";
when 1289 => read_data_o <= x"0064";
when 1290 => read_data_o <= x"0064";
when 1291 => read_data_o <= x"0064";
when 1292 => read_data_o <= x"0064";
when 1293 => read_data_o <= x"0064";
when 1294 => read_data_o <= x"0064";
when 1295 => read_data_o <= x"0064";
when 1296 => read_data_o <= x"0064";
when 1297 => read_data_o <= x"0064";
when 1298 => read_data_o <= x"0064";
when 1299 => read_data_o <= x"0064";
when 1300 => read_data_o <= x"0064";
when 1301 => read_data_o <= x"0064";
when 1302 => read_data_o <= x"0064";
when 1303 => read_data_o <= x"0064";
when 1304 => read_data_o <= x"0064";
when 1305 => read_data_o <= x"0064";
when 1306 => read_data_o <= x"0064";
when 1307 => read_data_o <= x"0064";
when 1308 => read_data_o <= x"0064";
when 1309 => read_data_o <= x"0064";
when 1310 => read_data_o <= x"0064";
when 1311 => read_data_o <= x"0064";
when 1312 => read_data_o <= x"0064";
when 1313 => read_data_o <= x"0064";
when 1314 => read_data_o <= x"0064";
when 1315 => read_data_o <= x"0064";
when 1316 => read_data_o <= x"0064";
when 1317 => read_data_o <= x"0064";
when 1318 => read_data_o <= x"0064";
when 1319 => read_data_o <= x"0064";
when 1320 => read_data_o <= x"0064";
when 1321 => read_data_o <= x"0064";
when 1322 => read_data_o <= x"0064";
when 1323 => read_data_o <= x"0064";
when 1324 => read_data_o <= x"0064";
when 1325 => read_data_o <= x"0064";
when 1326 => read_data_o <= x"0064";
when 1327 => read_data_o <= x"0064";
when 1328 => read_data_o <= x"0064";
when 1329 => read_data_o <= x"0064";
when 1330 => read_data_o <= x"0064";
when 1331 => read_data_o <= x"0064";
when 1332 => read_data_o <= x"0064";
when 1333 => read_data_o <= x"0064";
when 1334 => read_data_o <= x"0064";
when 1335 => read_data_o <= x"0064";
when 1336 => read_data_o <= x"0064";
when 1337 => read_data_o <= x"0064";
when 1338 => read_data_o <= x"0064";
when 1339 => read_data_o <= x"0064";
when 1340 => read_data_o <= x"0064";
when 1341 => read_data_o <= x"0064";
when 1342 => read_data_o <= x"0064";
when 1343 => read_data_o <= x"0064";
when 1344 => read_data_o <= x"0064";
when 1345 => read_data_o <= x"0064";
when 1346 => read_data_o <= x"0064";
when 1347 => read_data_o <= x"0064";
when 1348 => read_data_o <= x"0064";
when 1349 => read_data_o <= x"0064";
when 1350 => read_data_o <= x"0064";
when 1351 => read_data_o <= x"0064";
when 1352 => read_data_o <= x"0064";
when 1353 => read_data_o <= x"0064";
when 1354 => read_data_o <= x"0064";
when 1355 => read_data_o <= x"0064";
when 1356 => read_data_o <= x"0064";
when 1357 => read_data_o <= x"0064";
when 1358 => read_data_o <= x"0064";
when 1359 => read_data_o <= x"0064";
when 1360 => read_data_o <= x"0064";
when 1361 => read_data_o <= x"0064";
when 1362 => read_data_o <= x"0064";
when 1363 => read_data_o <= x"0064";
when 1364 => read_data_o <= x"0064";
when 1365 => read_data_o <= x"0064";
when 1366 => read_data_o <= x"0064";
when 1367 => read_data_o <= x"0064";
when 1368 => read_data_o <= x"0064";
when 1369 => read_data_o <= x"0064";
when 1370 => read_data_o <= x"0064";
when 1371 => read_data_o <= x"0064";
when 1372 => read_data_o <= x"0064";
when 1373 => read_data_o <= x"0064";
when 1374 => read_data_o <= x"0064";
when 1375 => read_data_o <= x"0064";
when 1376 => read_data_o <= x"0064";
when 1377 => read_data_o <= x"0064";
when 1378 => read_data_o <= x"0064";
when 1379 => read_data_o <= x"0064";
when 1380 => read_data_o <= x"0064";
when 1381 => read_data_o <= x"0064";
when 1382 => read_data_o <= x"0064";
when 1383 => read_data_o <= x"0064";
when 1384 => read_data_o <= x"0064";
when 1385 => read_data_o <= x"0064";
when 1386 => read_data_o <= x"0064";
when 1387 => read_data_o <= x"0064";
when 1388 => read_data_o <= x"0064";
when 1389 => read_data_o <= x"0064";
when 1390 => read_data_o <= x"0064";
when 1391 => read_data_o <= x"0064";
when 1392 => read_data_o <= x"0064";
when 1393 => read_data_o <= x"0064";
when 1394 => read_data_o <= x"0064";
when 1395 => read_data_o <= x"0064";
when 1396 => read_data_o <= x"0064";
when 1397 => read_data_o <= x"0064";
when 1398 => read_data_o <= x"0064";
when 1399 => read_data_o <= x"0064";
when 1400 => read_data_o <= x"0064";
when 1401 => read_data_o <= x"0064";
when 1402 => read_data_o <= x"0064";
when 1403 => read_data_o <= x"0064";
when 1404 => read_data_o <= x"0064";
when 1405 => read_data_o <= x"0064";
when 1406 => read_data_o <= x"0064";
when 1407 => read_data_o <= x"0064";
when 1408 => read_data_o <= x"0064";
when 1409 => read_data_o <= x"0064";
when 1410 => read_data_o <= x"0064";
when 1411 => read_data_o <= x"0064";
when 1412 => read_data_o <= x"0064";
when 1413 => read_data_o <= x"0064";
when 1414 => read_data_o <= x"0064";
when 1415 => read_data_o <= x"0064";
when 1416 => read_data_o <= x"0064";
when 1417 => read_data_o <= x"0064";
when 1418 => read_data_o <= x"0064";
when 1419 => read_data_o <= x"0064";
when 1420 => read_data_o <= x"0064";
when 1421 => read_data_o <= x"0064";
when 1422 => read_data_o <= x"0064";
when 1423 => read_data_o <= x"0064";
when 1424 => read_data_o <= x"0064";
when 1425 => read_data_o <= x"0064";
when 1426 => read_data_o <= x"0064";
when 1427 => read_data_o <= x"0064";
when 1428 => read_data_o <= x"0064";
when 1429 => read_data_o <= x"0064";
when 1430 => read_data_o <= x"0064";
when 1431 => read_data_o <= x"0064";
when 1432 => read_data_o <= x"0064";
when 1433 => read_data_o <= x"0064";
when 1434 => read_data_o <= x"0064";
when 1435 => read_data_o <= x"0064";
when 1436 => read_data_o <= x"0064";
when 1437 => read_data_o <= x"0064";
when 1438 => read_data_o <= x"0064";
when 1439 => read_data_o <= x"0064";
when 1440 => read_data_o <= x"0064";
when 1441 => read_data_o <= x"0064";
when 1442 => read_data_o <= x"0064";
when 1443 => read_data_o <= x"0064";
when 1444 => read_data_o <= x"0064";
when 1445 => read_data_o <= x"0064";
when 1446 => read_data_o <= x"0064";
when 1447 => read_data_o <= x"0064";
when 1448 => read_data_o <= x"0064";
when 1449 => read_data_o <= x"0064";
when 1450 => read_data_o <= x"0064";
when 1451 => read_data_o <= x"0064";
when 1452 => read_data_o <= x"0064";
when 1453 => read_data_o <= x"0064";
when 1454 => read_data_o <= x"0064";
when 1455 => read_data_o <= x"0064";
when 1456 => read_data_o <= x"0064";
when 1457 => read_data_o <= x"0064";
when 1458 => read_data_o <= x"0064";
when 1459 => read_data_o <= x"0064";
when 1460 => read_data_o <= x"0064";
when 1461 => read_data_o <= x"0064";
when 1462 => read_data_o <= x"0064";
when 1463 => read_data_o <= x"0064";
when 1464 => read_data_o <= x"0064";
when 1465 => read_data_o <= x"0064";
when 1466 => read_data_o <= x"0064";
when 1467 => read_data_o <= x"0064";
when 1468 => read_data_o <= x"0064";
when 1469 => read_data_o <= x"0064";
when 1470 => read_data_o <= x"0064";
when 1471 => read_data_o <= x"0064";
when 1472 => read_data_o <= x"0064";
when 1473 => read_data_o <= x"0064";
when 1474 => read_data_o <= x"0064";
when 1475 => read_data_o <= x"0064";
when 1476 => read_data_o <= x"0064";
when 1477 => read_data_o <= x"0064";
when 1478 => read_data_o <= x"0064";
when 1479 => read_data_o <= x"0064";
when 1480 => read_data_o <= x"0064";
when 1481 => read_data_o <= x"0064";
when 1482 => read_data_o <= x"0064";
when 1483 => read_data_o <= x"0064";
when 1484 => read_data_o <= x"0064";
when 1485 => read_data_o <= x"0064";
when 1486 => read_data_o <= x"0064";
when 1487 => read_data_o <= x"0064";
when 1488 => read_data_o <= x"0064";
when 1489 => read_data_o <= x"0064";
when 1490 => read_data_o <= x"0064";
when 1491 => read_data_o <= x"0064";
when 1492 => read_data_o <= x"0064";
when 1493 => read_data_o <= x"0064";
when 1494 => read_data_o <= x"0064";
when 1495 => read_data_o <= x"0064";
when 1496 => read_data_o <= x"0064";
when 1497 => read_data_o <= x"0064";
when 1498 => read_data_o <= x"0064";
when 1499 => read_data_o <= x"0064";
when 1500 => read_data_o <= x"0064";
when 1501 => read_data_o <= x"0064";
when 1502 => read_data_o <= x"0064";
when 1503 => read_data_o <= x"0064";
when 1504 => read_data_o <= x"0064";
when 1505 => read_data_o <= x"0064";
when 1506 => read_data_o <= x"0064";
when 1507 => read_data_o <= x"0064";
when 1508 => read_data_o <= x"0064";
when 1509 => read_data_o <= x"0064";
when 1510 => read_data_o <= x"0064";
when 1511 => read_data_o <= x"0064";
when 1512 => read_data_o <= x"0064";
when 1513 => read_data_o <= x"0064";
when 1514 => read_data_o <= x"0064";
when 1515 => read_data_o <= x"0064";
when 1516 => read_data_o <= x"0064";
when 1517 => read_data_o <= x"0064";
when 1518 => read_data_o <= x"0064";
when 1519 => read_data_o <= x"0064";
when 1520 => read_data_o <= x"0064";
when 1521 => read_data_o <= x"0064";
when 1522 => read_data_o <= x"0064";
when 1523 => read_data_o <= x"0064";
when 1524 => read_data_o <= x"0064";
when 1525 => read_data_o <= x"0064";
when 1526 => read_data_o <= x"0064";
when 1527 => read_data_o <= x"0064";
when 1528 => read_data_o <= x"0064";
when 1529 => read_data_o <= x"0064";
when 1530 => read_data_o <= x"0064";
when 1531 => read_data_o <= x"0064";
when 1532 => read_data_o <= x"0064";
when 1533 => read_data_o <= x"0064";
when 1534 => read_data_o <= x"0064";
when 1535 => read_data_o <= x"0064";
when 1536 => read_data_o <= x"0064";
when 1537 => read_data_o <= x"0064";
when 1538 => read_data_o <= x"0064";
when 1539 => read_data_o <= x"0064";
when 1540 => read_data_o <= x"0064";
when 1541 => read_data_o <= x"0064";
when 1542 => read_data_o <= x"0064";
when 1543 => read_data_o <= x"0064";
when 1544 => read_data_o <= x"0064";
when 1545 => read_data_o <= x"0064";
when 1546 => read_data_o <= x"0064";
when 1547 => read_data_o <= x"0064";
when 1548 => read_data_o <= x"0064";
when 1549 => read_data_o <= x"0064";
when 1550 => read_data_o <= x"0064";
when 1551 => read_data_o <= x"0064";
when 1552 => read_data_o <= x"0064";
when 1553 => read_data_o <= x"0064";
when 1554 => read_data_o <= x"0064";
when 1555 => read_data_o <= x"0064";
when 1556 => read_data_o <= x"0064";
when 1557 => read_data_o <= x"0064";
when 1558 => read_data_o <= x"0064";
when 1559 => read_data_o <= x"0064";
when 1560 => read_data_o <= x"0064";
when 1561 => read_data_o <= x"0064";
when 1562 => read_data_o <= x"0064";
when 1563 => read_data_o <= x"0064";
when 1564 => read_data_o <= x"0064";
when 1565 => read_data_o <= x"0064";
when 1566 => read_data_o <= x"0064";
when 1567 => read_data_o <= x"0064";
when 1568 => read_data_o <= x"0064";
when 1569 => read_data_o <= x"0064";
when 1570 => read_data_o <= x"0064";
when 1571 => read_data_o <= x"0064";
when 1572 => read_data_o <= x"0064";
when 1573 => read_data_o <= x"0064";
when 1574 => read_data_o <= x"0064";
when 1575 => read_data_o <= x"0064";
when 1576 => read_data_o <= x"0064";
when 1577 => read_data_o <= x"0064";
when 1578 => read_data_o <= x"0064";
when 1579 => read_data_o <= x"0064";
when 1580 => read_data_o <= x"0064";
when 1581 => read_data_o <= x"0064";
when 1582 => read_data_o <= x"0064";
when 1583 => read_data_o <= x"0064";
when 1584 => read_data_o <= x"0064";
when 1585 => read_data_o <= x"0064";
when 1586 => read_data_o <= x"0064";
when 1587 => read_data_o <= x"0064";
when 1588 => read_data_o <= x"0064";
when 1589 => read_data_o <= x"0064";
when 1590 => read_data_o <= x"0064";
when 1591 => read_data_o <= x"0064";
when 1592 => read_data_o <= x"0064";
when 1593 => read_data_o <= x"0064";
when 1594 => read_data_o <= x"0064";
when 1595 => read_data_o <= x"0064";
when 1596 => read_data_o <= x"0064";
when 1597 => read_data_o <= x"0064";
when 1598 => read_data_o <= x"0064";
when 1599 => read_data_o <= x"0064";
when 1600 => read_data_o <= x"0064";
when 1601 => read_data_o <= x"0064";
when 1602 => read_data_o <= x"0064";
when 1603 => read_data_o <= x"0064";
when 1604 => read_data_o <= x"0064";
when 1605 => read_data_o <= x"0064";
when 1606 => read_data_o <= x"0064";
when 1607 => read_data_o <= x"0064";
when 1608 => read_data_o <= x"0064";
when 1609 => read_data_o <= x"0064";
when 1610 => read_data_o <= x"0064";
when 1611 => read_data_o <= x"0064";
when 1612 => read_data_o <= x"2000";
when 1613 => read_data_o <= x"2000";
when 1614 => read_data_o <= x"2000";
when 1615 => read_data_o <= x"2000";
when 1616 => read_data_o <= x"2000";
when 1617 => read_data_o <= x"2405";
when 1618 => read_data_o <= x"7064";
when 1619 => read_data_o <= x"3064";
when 1620 => read_data_o <= x"3064";
when 1621 => read_data_o <= x"3064";
when 1622 => read_data_o <= x"3064";
when 1623 => read_data_o <= x"3064";
when 1624 => read_data_o <= x"3064";
when 1625 => read_data_o <= x"3064";
when 1626 => read_data_o <= x"3064";
when 1627 => read_data_o <= x"3064";
when 1628 => read_data_o <= x"3064";
when 1629 => read_data_o <= x"3064";
when 1630 => read_data_o <= x"3064";
when 1631 => read_data_o <= x"3064";
when 1632 => read_data_o <= x"3064";
when 1633 => read_data_o <= x"3064";
when 1634 => read_data_o <= x"3064";
when 1635 => read_data_o <= x"3064";
when 1636 => read_data_o <= x"3064";
when 1637 => read_data_o <= x"3064";
when 1638 => read_data_o <= x"3064";
when 1639 => read_data_o <= x"3064";
when 1640 => read_data_o <= x"3064";
when 1641 => read_data_o <= x"3064";
when 1642 => read_data_o <= x"3064";
when 1643 => read_data_o <= x"3064";
when 1644 => read_data_o <= x"3064";
when 1645 => read_data_o <= x"3064";
when 1646 => read_data_o <= x"3064";
when 1647 => read_data_o <= x"3064";
when 1648 => read_data_o <= x"3064";
when 1649 => read_data_o <= x"3064";
when 1650 => read_data_o <= x"3064";
when 1651 => read_data_o <= x"3064";
when 1652 => read_data_o <= x"3064";
when 1653 => read_data_o <= x"3064";
when 1654 => read_data_o <= x"3064";
when 1655 => read_data_o <= x"3064";
when 1656 => read_data_o <= x"3064";
when 1657 => read_data_o <= x"3064";
when 1658 => read_data_o <= x"3064";
when 1659 => read_data_o <= x"3064";
when 1660 => read_data_o <= x"3064";
when 1661 => read_data_o <= x"3064";
when 1662 => read_data_o <= x"3064";
when 1663 => read_data_o <= x"3064";
when 1664 => read_data_o <= x"3064";
when 1665 => read_data_o <= x"3064";
when 1666 => read_data_o <= x"3064";
when 1667 => read_data_o <= x"3064";
when 1668 => read_data_o <= x"3064";
when 1669 => read_data_o <= x"3064";
when 1670 => read_data_o <= x"3064";
when 1671 => read_data_o <= x"3064";
when 1672 => read_data_o <= x"3064";
when 1673 => read_data_o <= x"3064";
when 1674 => read_data_o <= x"3064";
when 1675 => read_data_o <= x"3064";
when 1676 => read_data_o <= x"3064";
when 1677 => read_data_o <= x"3064";
when 1678 => read_data_o <= x"3064";
when 1679 => read_data_o <= x"3064";
when 1680 => read_data_o <= x"3064";
when 1681 => read_data_o <= x"3064";
when 1682 => read_data_o <= x"3064";
when 1683 => read_data_o <= x"3064";
when 1684 => read_data_o <= x"3064";
when 1685 => read_data_o <= x"3064";
when 1686 => read_data_o <= x"3064";
when 1687 => read_data_o <= x"3064";
when 1688 => read_data_o <= x"3064";
when 1689 => read_data_o <= x"3064";
when 1690 => read_data_o <= x"3064";
when 1691 => read_data_o <= x"3064";
when 1692 => read_data_o <= x"3064";
when 1693 => read_data_o <= x"3064";
when 1694 => read_data_o <= x"3064";
when 1695 => read_data_o <= x"3064";
when 1696 => read_data_o <= x"3064";
when 1697 => read_data_o <= x"3064";
when 1698 => read_data_o <= x"3064";
when 1699 => read_data_o <= x"3064";
when 1700 => read_data_o <= x"3064";
when 1701 => read_data_o <= x"3064";
when 1702 => read_data_o <= x"3064";
when 1703 => read_data_o <= x"3064";
when 1704 => read_data_o <= x"3064";
when 1705 => read_data_o <= x"3064";
when 1706 => read_data_o <= x"3064";
when 1707 => read_data_o <= x"3064";
when 1708 => read_data_o <= x"3064";
when 1709 => read_data_o <= x"3064";
when 1710 => read_data_o <= x"3064";
when 1711 => read_data_o <= x"3064";
when 1712 => read_data_o <= x"3064";
when 1713 => read_data_o <= x"3064";
when 1714 => read_data_o <= x"3064";
when 1715 => read_data_o <= x"3064";
when 1716 => read_data_o <= x"3064";
when 1717 => read_data_o <= x"3064";
when 1718 => read_data_o <= x"3064";
when 1719 => read_data_o <= x"3064";
when 1720 => read_data_o <= x"3064";
when 1721 => read_data_o <= x"3064";
when 1722 => read_data_o <= x"3064";
when 1723 => read_data_o <= x"3064";
when 1724 => read_data_o <= x"3064";
when 1725 => read_data_o <= x"3064";
when 1726 => read_data_o <= x"3064";
when 1727 => read_data_o <= x"3064";
when 1728 => read_data_o <= x"3064";
when 1729 => read_data_o <= x"3064";
when 1730 => read_data_o <= x"3064";
when 1731 => read_data_o <= x"3064";
when 1732 => read_data_o <= x"3064";
when 1733 => read_data_o <= x"3064";
when 1734 => read_data_o <= x"3064";
when 1735 => read_data_o <= x"3064";
when 1736 => read_data_o <= x"3064";
when 1737 => read_data_o <= x"3064";
when 1738 => read_data_o <= x"3064";
when 1739 => read_data_o <= x"3064";
when 1740 => read_data_o <= x"3064";
when 1741 => read_data_o <= x"3064";
when 1742 => read_data_o <= x"3064";
when 1743 => read_data_o <= x"3064";
when 1744 => read_data_o <= x"3064";
when 1745 => read_data_o <= x"3064";
when 1746 => read_data_o <= x"3064";
when 1747 => read_data_o <= x"3064";
when 1748 => read_data_o <= x"3064";
when 1749 => read_data_o <= x"3064";
when 1750 => read_data_o <= x"3064";
when 1751 => read_data_o <= x"3064";
when 1752 => read_data_o <= x"3064";
when 1753 => read_data_o <= x"3064";
when 1754 => read_data_o <= x"3064";
when 1755 => read_data_o <= x"3064";
when 1756 => read_data_o <= x"3064";
when 1757 => read_data_o <= x"3064";
when 1758 => read_data_o <= x"3064";
when 1759 => read_data_o <= x"3064";
when 1760 => read_data_o <= x"3064";
when 1761 => read_data_o <= x"3064";
when 1762 => read_data_o <= x"3064";
when 1763 => read_data_o <= x"3064";
when 1764 => read_data_o <= x"3064";
when 1765 => read_data_o <= x"3064";
when 1766 => read_data_o <= x"3064";
when 1767 => read_data_o <= x"3064";
when 1768 => read_data_o <= x"3064";
when 1769 => read_data_o <= x"3064";
when 1770 => read_data_o <= x"3064";
when 1771 => read_data_o <= x"3064";
when 1772 => read_data_o <= x"3064";
when 1773 => read_data_o <= x"3064";
when 1774 => read_data_o <= x"3064";
when 1775 => read_data_o <= x"3064";
when 1776 => read_data_o <= x"3064";
when 1777 => read_data_o <= x"3064";
when 1778 => read_data_o <= x"3064";
when 1779 => read_data_o <= x"3064";
when 1780 => read_data_o <= x"3064";
when 1781 => read_data_o <= x"3064";
when 1782 => read_data_o <= x"3064";
when 1783 => read_data_o <= x"3064";
when 1784 => read_data_o <= x"3064";
when 1785 => read_data_o <= x"3064";
when 1786 => read_data_o <= x"3064";
when 1787 => read_data_o <= x"3064";
when 1788 => read_data_o <= x"3064";
when 1789 => read_data_o <= x"3064";
when 1790 => read_data_o <= x"3064";
when 1791 => read_data_o <= x"3064";
when 1792 => read_data_o <= x"3064";
when 1793 => read_data_o <= x"3064";
when 1794 => read_data_o <= x"3064";
when 1795 => read_data_o <= x"3064";
when 1796 => read_data_o <= x"3064";
when 1797 => read_data_o <= x"3064";
when 1798 => read_data_o <= x"3064";
when 1799 => read_data_o <= x"3064";
when 1800 => read_data_o <= x"3064";
when 1801 => read_data_o <= x"3064";
when 1802 => read_data_o <= x"3064";
when 1803 => read_data_o <= x"3064";
when 1804 => read_data_o <= x"3064";
when 1805 => read_data_o <= x"3064";
when 1806 => read_data_o <= x"3064";
when 1807 => read_data_o <= x"3064";
when 1808 => read_data_o <= x"3064";
when 1809 => read_data_o <= x"3064";
when 1810 => read_data_o <= x"3064";
when 1811 => read_data_o <= x"3064";
when 1812 => read_data_o <= x"3064";
when 1813 => read_data_o <= x"3064";
when 1814 => read_data_o <= x"3064";
when 1815 => read_data_o <= x"3064";
when 1816 => read_data_o <= x"3064";
when 1817 => read_data_o <= x"3064";
when 1818 => read_data_o <= x"3064";
when 1819 => read_data_o <= x"3064";
when 1820 => read_data_o <= x"3064";
when 1821 => read_data_o <= x"3064";
when 1822 => read_data_o <= x"3064";
when 1823 => read_data_o <= x"3064";
when 1824 => read_data_o <= x"3064";
when 1825 => read_data_o <= x"3064";
when 1826 => read_data_o <= x"3064";
when 1827 => read_data_o <= x"3064";
when 1828 => read_data_o <= x"3064";
when 1829 => read_data_o <= x"3064";
when 1830 => read_data_o <= x"3064";
when 1831 => read_data_o <= x"3064";
when 1832 => read_data_o <= x"3064";
when 1833 => read_data_o <= x"3064";
when 1834 => read_data_o <= x"3064";
when 1835 => read_data_o <= x"3064";
when 1836 => read_data_o <= x"3064";
when 1837 => read_data_o <= x"3064";
when 1838 => read_data_o <= x"3064";
when 1839 => read_data_o <= x"3064";
when 1840 => read_data_o <= x"3064";
when 1841 => read_data_o <= x"3064";
when 1842 => read_data_o <= x"3064";
when 1843 => read_data_o <= x"3064";
when 1844 => read_data_o <= x"3064";
when 1845 => read_data_o <= x"3064";
when 1846 => read_data_o <= x"3064";
when 1847 => read_data_o <= x"3064";
when 1848 => read_data_o <= x"3064";
when 1849 => read_data_o <= x"3064";
when 1850 => read_data_o <= x"3064";
when 1851 => read_data_o <= x"3064";
when 1852 => read_data_o <= x"3064";
when 1853 => read_data_o <= x"3064";
when 1854 => read_data_o <= x"3064";
when 1855 => read_data_o <= x"3064";
when 1856 => read_data_o <= x"3064";
when 1857 => read_data_o <= x"3064";
when 1858 => read_data_o <= x"3064";
when 1859 => read_data_o <= x"3064";
when 1860 => read_data_o <= x"3064";
when 1861 => read_data_o <= x"3064";
when 1862 => read_data_o <= x"3064";
when 1863 => read_data_o <= x"3064";
when 1864 => read_data_o <= x"3064";
when 1865 => read_data_o <= x"3064";
when 1866 => read_data_o <= x"3064";
when 1867 => read_data_o <= x"3064";
when 1868 => read_data_o <= x"3064";
when 1869 => read_data_o <= x"3064";
when 1870 => read_data_o <= x"3064";
when 1871 => read_data_o <= x"3064";
when 1872 => read_data_o <= x"3064";
when 1873 => read_data_o <= x"3064";
when 1874 => read_data_o <= x"3064";
when 1875 => read_data_o <= x"3064";
when 1876 => read_data_o <= x"3064";
when 1877 => read_data_o <= x"3064";
when 1878 => read_data_o <= x"3064";
when 1879 => read_data_o <= x"3064";
when 1880 => read_data_o <= x"3064";
when 1881 => read_data_o <= x"3064";
when 1882 => read_data_o <= x"3064";
when 1883 => read_data_o <= x"3064";
when 1884 => read_data_o <= x"3064";
when 1885 => read_data_o <= x"3064";
when 1886 => read_data_o <= x"3064";
when 1887 => read_data_o <= x"3064";
when 1888 => read_data_o <= x"3064";
when 1889 => read_data_o <= x"3064";
when 1890 => read_data_o <= x"3064";
when 1891 => read_data_o <= x"3064";
when 1892 => read_data_o <= x"3064";
when 1893 => read_data_o <= x"3064";
when 1894 => read_data_o <= x"3064";
when 1895 => read_data_o <= x"3064";
when 1896 => read_data_o <= x"3064";
when 1897 => read_data_o <= x"3064";
when 1898 => read_data_o <= x"3064";
when 1899 => read_data_o <= x"3064";
when 1900 => read_data_o <= x"3064";
when 1901 => read_data_o <= x"3064";
when 1902 => read_data_o <= x"3064";
when 1903 => read_data_o <= x"3064";
when 1904 => read_data_o <= x"3064";
when 1905 => read_data_o <= x"3064";
when 1906 => read_data_o <= x"3064";
when 1907 => read_data_o <= x"3064";
when 1908 => read_data_o <= x"3064";
when 1909 => read_data_o <= x"3064";
when 1910 => read_data_o <= x"3064";
when 1911 => read_data_o <= x"3064";
when 1912 => read_data_o <= x"3064";
when 1913 => read_data_o <= x"3064";
when 1914 => read_data_o <= x"3064";
when 1915 => read_data_o <= x"3064";
when 1916 => read_data_o <= x"3064";
when 1917 => read_data_o <= x"3064";
when 1918 => read_data_o <= x"3064";
when 1919 => read_data_o <= x"3064";
when 1920 => read_data_o <= x"3064";
when 1921 => read_data_o <= x"3064";
when 1922 => read_data_o <= x"3064";
when 1923 => read_data_o <= x"3064";
when 1924 => read_data_o <= x"3064";
when 1925 => read_data_o <= x"3064";
when 1926 => read_data_o <= x"3064";
when 1927 => read_data_o <= x"3064";
when 1928 => read_data_o <= x"3064";
when 1929 => read_data_o <= x"3064";
when 1930 => read_data_o <= x"3064";
when 1931 => read_data_o <= x"3064";
when 1932 => read_data_o <= x"3064";
when 1933 => read_data_o <= x"3064";
when 1934 => read_data_o <= x"3064";
when 1935 => read_data_o <= x"3064";
when 1936 => read_data_o <= x"3064";
when 1937 => read_data_o <= x"3064";
when 1938 => read_data_o <= x"3064";
when 1939 => read_data_o <= x"3064";
when 1940 => read_data_o <= x"3064";
when 1941 => read_data_o <= x"3064";
when 1942 => read_data_o <= x"3064";
when 1943 => read_data_o <= x"3064";
when 1944 => read_data_o <= x"3064";
when 1945 => read_data_o <= x"3064";
when 1946 => read_data_o <= x"3064";
when 1947 => read_data_o <= x"3064";
when 1948 => read_data_o <= x"3064";
when 1949 => read_data_o <= x"3064";
when 1950 => read_data_o <= x"3064";
when 1951 => read_data_o <= x"3064";
when 1952 => read_data_o <= x"3064";
when 1953 => read_data_o <= x"3064";
when 1954 => read_data_o <= x"3064";
when 1955 => read_data_o <= x"3064";
when 1956 => read_data_o <= x"3064";
when 1957 => read_data_o <= x"3064";
when 1958 => read_data_o <= x"3064";
when 1959 => read_data_o <= x"3064";
when 1960 => read_data_o <= x"3064";
when 1961 => read_data_o <= x"3064";
when 1962 => read_data_o <= x"3064";
when 1963 => read_data_o <= x"3064";
when 1964 => read_data_o <= x"3064";
when 1965 => read_data_o <= x"3064";
when 1966 => read_data_o <= x"3064";
when 1967 => read_data_o <= x"3064";
when 1968 => read_data_o <= x"3064";
when 1969 => read_data_o <= x"3064";
when 1970 => read_data_o <= x"3064";
when 1971 => read_data_o <= x"3064";
when 1972 => read_data_o <= x"3064";
when 1973 => read_data_o <= x"3064";
when 1974 => read_data_o <= x"3064";
when 1975 => read_data_o <= x"3064";
when 1976 => read_data_o <= x"3064";
when 1977 => read_data_o <= x"3064";
when 1978 => read_data_o <= x"3064";
when 1979 => read_data_o <= x"3064";
when 1980 => read_data_o <= x"3064";
when 1981 => read_data_o <= x"3064";
when 1982 => read_data_o <= x"3064";
when 1983 => read_data_o <= x"3064";
when 1984 => read_data_o <= x"3064";
when 1985 => read_data_o <= x"3064";
when 1986 => read_data_o <= x"3064";
when 1987 => read_data_o <= x"3064";
when 1988 => read_data_o <= x"3064";
when 1989 => read_data_o <= x"3064";
when 1990 => read_data_o <= x"3064";
when 1991 => read_data_o <= x"3064";
when 1992 => read_data_o <= x"3064";
when 1993 => read_data_o <= x"3064";
when 1994 => read_data_o <= x"3064";
when 1995 => read_data_o <= x"3064";
when 1996 => read_data_o <= x"3064";
when 1997 => read_data_o <= x"3064";
when 1998 => read_data_o <= x"3064";
when 1999 => read_data_o <= x"3064";
when 2000 => read_data_o <= x"3064";
when 2001 => read_data_o <= x"3064";
when 2002 => read_data_o <= x"3064";
when 2003 => read_data_o <= x"3064";
when 2004 => read_data_o <= x"3064";
when 2005 => read_data_o <= x"3064";
when 2006 => read_data_o <= x"3064";
when 2007 => read_data_o <= x"3064";
when 2008 => read_data_o <= x"3064";
when 2009 => read_data_o <= x"3064";
when 2010 => read_data_o <= x"3064";
when 2011 => read_data_o <= x"3064";
when 2012 => read_data_o <= x"3064";
when 2013 => read_data_o <= x"3064";
when 2014 => read_data_o <= x"3064";
when 2015 => read_data_o <= x"3064";
when 2016 => read_data_o <= x"3064";
when 2017 => read_data_o <= x"3064";
when 2018 => read_data_o <= x"3064";
when 2019 => read_data_o <= x"3064";
when 2020 => read_data_o <= x"3064";
when 2021 => read_data_o <= x"3064";
when 2022 => read_data_o <= x"3064";
when 2023 => read_data_o <= x"3064";
when 2024 => read_data_o <= x"3064";
when 2025 => read_data_o <= x"3064";
when 2026 => read_data_o <= x"3064";
when 2027 => read_data_o <= x"3064";
when 2028 => read_data_o <= x"3064";
when 2029 => read_data_o <= x"3064";
when 2030 => read_data_o <= x"3064";
when 2031 => read_data_o <= x"3064";
when 2032 => read_data_o <= x"3064";
when 2033 => read_data_o <= x"3064";
when 2034 => read_data_o <= x"3064";
when 2035 => read_data_o <= x"3064";
when 2036 => read_data_o <= x"3064";
when 2037 => read_data_o <= x"3064";
when 2038 => read_data_o <= x"3064";
when 2039 => read_data_o <= x"3064";
when 2040 => read_data_o <= x"3064";
when 2041 => read_data_o <= x"3064";
when 2042 => read_data_o <= x"3064";
when 2043 => read_data_o <= x"3064";
when 2044 => read_data_o <= x"3064";
when 2045 => read_data_o <= x"3064";
when 2046 => read_data_o <= x"3064";
when 2047 => read_data_o <= x"3064";
when 2048 => read_data_o <= x"3064";
when 2049 => read_data_o <= x"3064";
when 2050 => read_data_o <= x"3064";
when 2051 => read_data_o <= x"3064";
when 2052 => read_data_o <= x"3064";
when 2053 => read_data_o <= x"3064";
when 2054 => read_data_o <= x"3064";
when 2055 => read_data_o <= x"3064";
when 2056 => read_data_o <= x"3064";
when 2057 => read_data_o <= x"3064";
when 2058 => read_data_o <= x"3064";
when 2059 => read_data_o <= x"3064";
when 2060 => read_data_o <= x"3064";
when 2061 => read_data_o <= x"3064";
when 2062 => read_data_o <= x"3064";
when 2063 => read_data_o <= x"3064";
when 2064 => read_data_o <= x"3064";
when 2065 => read_data_o <= x"3064";
when 2066 => read_data_o <= x"3064";
when 2067 => read_data_o <= x"3064";
when 2068 => read_data_o <= x"3064";
when 2069 => read_data_o <= x"3064";
when 2070 => read_data_o <= x"3064";
when 2071 => read_data_o <= x"3064";
when 2072 => read_data_o <= x"3064";
when 2073 => read_data_o <= x"3064";
when 2074 => read_data_o <= x"3064";
when 2075 => read_data_o <= x"3064";
when 2076 => read_data_o <= x"3064";
when 2077 => read_data_o <= x"3064";
when 2078 => read_data_o <= x"3064";
when 2079 => read_data_o <= x"3064";
when 2080 => read_data_o <= x"3064";
when 2081 => read_data_o <= x"3064";
when 2082 => read_data_o <= x"3064";
when 2083 => read_data_o <= x"3064";
when 2084 => read_data_o <= x"3064";
when 2085 => read_data_o <= x"3064";
when 2086 => read_data_o <= x"3064";
when 2087 => read_data_o <= x"3064";
when 2088 => read_data_o <= x"3064";
when 2089 => read_data_o <= x"3064";
when 2090 => read_data_o <= x"3064";
when 2091 => read_data_o <= x"3064";
when 2092 => read_data_o <= x"3064";
when 2093 => read_data_o <= x"3064";
when 2094 => read_data_o <= x"3064";
when 2095 => read_data_o <= x"3064";
when 2096 => read_data_o <= x"3064";
when 2097 => read_data_o <= x"3064";
when 2098 => read_data_o <= x"3064";
when 2099 => read_data_o <= x"3064";
when 2100 => read_data_o <= x"3064";
when 2101 => read_data_o <= x"3064";
when 2102 => read_data_o <= x"3064";
when 2103 => read_data_o <= x"3064";
when 2104 => read_data_o <= x"3064";
when 2105 => read_data_o <= x"3064";
when 2106 => read_data_o <= x"3064";
when 2107 => read_data_o <= x"3064";
when 2108 => read_data_o <= x"3064";
when 2109 => read_data_o <= x"3064";
when 2110 => read_data_o <= x"3064";
when 2111 => read_data_o <= x"3064";
when 2112 => read_data_o <= x"3064";
when 2113 => read_data_o <= x"3064";
when 2114 => read_data_o <= x"3064";
when 2115 => read_data_o <= x"3064";
when 2116 => read_data_o <= x"3064";
when 2117 => read_data_o <= x"3064";
when 2118 => read_data_o <= x"3064";
when 2119 => read_data_o <= x"3064";
when 2120 => read_data_o <= x"3064";
when 2121 => read_data_o <= x"3064";
when 2122 => read_data_o <= x"3064";
when 2123 => read_data_o <= x"3064";
when 2124 => read_data_o <= x"3064";
when 2125 => read_data_o <= x"3064";
when 2126 => read_data_o <= x"3064";
when 2127 => read_data_o <= x"3064";
when 2128 => read_data_o <= x"3064";
when 2129 => read_data_o <= x"3064";
when 2130 => read_data_o <= x"3064";
when 2131 => read_data_o <= x"3064";
when 2132 => read_data_o <= x"3064";
when 2133 => read_data_o <= x"3064";
when 2134 => read_data_o <= x"3064";
when 2135 => read_data_o <= x"3064";
when 2136 => read_data_o <= x"3064";
when 2137 => read_data_o <= x"3064";
when 2138 => read_data_o <= x"3064";
when 2139 => read_data_o <= x"3064";
when 2140 => read_data_o <= x"3064";
when 2141 => read_data_o <= x"3064";
when 2142 => read_data_o <= x"3064";
when 2143 => read_data_o <= x"3064";
when 2144 => read_data_o <= x"3064";
when 2145 => read_data_o <= x"3064";
when 2146 => read_data_o <= x"3064";
when 2147 => read_data_o <= x"3064";
when 2148 => read_data_o <= x"3064";
when 2149 => read_data_o <= x"3064";
when 2150 => read_data_o <= x"3064";
when 2151 => read_data_o <= x"3064";
when 2152 => read_data_o <= x"3064";
when 2153 => read_data_o <= x"3064";
when 2154 => read_data_o <= x"3064";
when 2155 => read_data_o <= x"3064";
when 2156 => read_data_o <= x"3064";
when 2157 => read_data_o <= x"3064";
when 2158 => read_data_o <= x"3064";
when 2159 => read_data_o <= x"3064";
when 2160 => read_data_o <= x"3064";
when 2161 => read_data_o <= x"3064";
when 2162 => read_data_o <= x"3064";
when 2163 => read_data_o <= x"3064";
when 2164 => read_data_o <= x"3064";
when 2165 => read_data_o <= x"3064";
when 2166 => read_data_o <= x"3064";
when 2167 => read_data_o <= x"3064";
when 2168 => read_data_o <= x"3064";
when 2169 => read_data_o <= x"3064";
when 2170 => read_data_o <= x"3064";
when 2171 => read_data_o <= x"3064";
when 2172 => read_data_o <= x"3064";
when 2173 => read_data_o <= x"3064";
when 2174 => read_data_o <= x"3064";
when 2175 => read_data_o <= x"3064";
when 2176 => read_data_o <= x"3064";
when 2177 => read_data_o <= x"3064";
when 2178 => read_data_o <= x"3064";
when 2179 => read_data_o <= x"3064";
when 2180 => read_data_o <= x"3064";
when 2181 => read_data_o <= x"3064";
when 2182 => read_data_o <= x"3064";
when 2183 => read_data_o <= x"3064";
when 2184 => read_data_o <= x"3064";
when 2185 => read_data_o <= x"3064";
when 2186 => read_data_o <= x"3064";
when 2187 => read_data_o <= x"3064";
when 2188 => read_data_o <= x"3064";
when 2189 => read_data_o <= x"3064";
when 2190 => read_data_o <= x"3064";
when 2191 => read_data_o <= x"3064";
when 2192 => read_data_o <= x"3064";
when 2193 => read_data_o <= x"3064";
when 2194 => read_data_o <= x"3064";
when 2195 => read_data_o <= x"3064";
when 2196 => read_data_o <= x"3064";
when 2197 => read_data_o <= x"3064";
when 2198 => read_data_o <= x"3064";
when 2199 => read_data_o <= x"3064";
when 2200 => read_data_o <= x"3064";
when 2201 => read_data_o <= x"3064";
when 2202 => read_data_o <= x"3064";
when 2203 => read_data_o <= x"3064";
when 2204 => read_data_o <= x"3064";
when 2205 => read_data_o <= x"3064";
when 2206 => read_data_o <= x"3064";
when 2207 => read_data_o <= x"3064";
when 2208 => read_data_o <= x"3064";
when 2209 => read_data_o <= x"3064";
when 2210 => read_data_o <= x"3064";
when 2211 => read_data_o <= x"3064";
when 2212 => read_data_o <= x"3064";
when 2213 => read_data_o <= x"3064";
when 2214 => read_data_o <= x"3064";
when 2215 => read_data_o <= x"3064";
when 2216 => read_data_o <= x"3064";
when 2217 => read_data_o <= x"3064";
when 2218 => read_data_o <= x"3064";
when 2219 => read_data_o <= x"3064";
when 2220 => read_data_o <= x"2000";
when 2221 => read_data_o <= x"2000";
when 2222 => read_data_o <= x"2000";
when 2223 => read_data_o <= x"2000";
when 2224 => read_data_o <= x"2000";
when 2225 => read_data_o <= x"b196";
when 2226 => read_data_o <= x"7064";
when 2227 => read_data_o <= x"02bc";
when 2228 => read_data_o <= x"a000";
when 2229 => read_data_o <= x"a000";
when 2230 => read_data_o <= x"a000";
when 2231 => read_data_o <= x"a000";
when 2232 => read_data_o <= x"a000";
when 2233 => read_data_o <= x"a000";
when 2234 => read_data_o <= x"a000";
when 2235 => read_data_o <= x"a000";
when 2236 => read_data_o <= x"a000";
when 2237 => read_data_o <= x"a000";
when 2238 => read_data_o <= x"a000";
when 2239 => read_data_o <= x"a000";
when 2240 => read_data_o <= x"a000";
when 2241 => read_data_o <= x"a000";
when 2242 => read_data_o <= x"a000";
when 2243 => read_data_o <= x"a000";
when 2244 => read_data_o <= x"a000";
when 2245 => read_data_o <= x"a000";
when 2246 => read_data_o <= x"a000";
when 2247 => read_data_o <= x"a000";
when 2248 => read_data_o <= x"a000";
when 2249 => read_data_o <= x"a000";
when 2250 => read_data_o <= x"a000";
when 2251 => read_data_o <= x"a000";
when 2252 => read_data_o <= x"2404";
when 2253 => read_data_o <= x"0000";
when 2254 => read_data_o <= x"2000";
when 2255 => read_data_o <= x"2000";
when 2256 => read_data_o <= x"2000";
when 2257 => read_data_o <= x"2000";
when 2258 => read_data_o <= x"2000";
when 2259 => read_data_o <= x"2000";
when 2260 => read_data_o <= x"2000";
when 2261 => read_data_o <= x"2000";
when 2262 => read_data_o <= x"2000";
when 2263 => read_data_o <= x"2000";
when 2264 => read_data_o <= x"2000";
when 2265 => read_data_o <= x"2000";
when 2266 => read_data_o <= x"2000";
when 2267 => read_data_o <= x"2000";
when 2268 => read_data_o <= x"2000";
when 2269 => read_data_o <= x"2000";
when 2270 => read_data_o <= x"2000";
when 2271 => read_data_o <= x"2000";
when 2272 => read_data_o <= x"2000";
when 2273 => read_data_o <= x"2000";
when 2274 => read_data_o <= x"2000";
when 2275 => read_data_o <= x"2000";
when 2276 => read_data_o <= x"2000";
when 2277 => read_data_o <= x"2000";
when 2278 => read_data_o <= x"2000";
when 2279 => read_data_o <= x"2000";
when 2280 => read_data_o <= x"2000";
when 2281 => read_data_o <= x"2000";
when 2282 => read_data_o <= x"2000";
when 2283 => read_data_o <= x"2000";
when 2284 => read_data_o <= x"2000";
when 2285 => read_data_o <= x"2000";
when 2286 => read_data_o <= x"2000";
when 2287 => read_data_o <= x"2000";
when 2288 => read_data_o <= x"2000";
when 2289 => read_data_o <= x"2000";
when 2290 => read_data_o <= x"2000";
when 2291 => read_data_o <= x"2000";
when 2292 => read_data_o <= x"2000";
when 2293 => read_data_o <= x"2000";
when 2294 => read_data_o <= x"2000";
when 2295 => read_data_o <= x"2000";
when 2296 => read_data_o <= x"2000";
when 2297 => read_data_o <= x"2000";
when 2298 => read_data_o <= x"2000";
when 2299 => read_data_o <= x"2000";
when 2300 => read_data_o <= x"2000";
when 2301 => read_data_o <= x"2000";
when 2302 => read_data_o <= x"2000";
when 2303 => read_data_o <= x"2000";
when 2304 => read_data_o <= x"2000";
when 2305 => read_data_o <= x"2000";
when 2306 => read_data_o <= x"2000";
when 2307 => read_data_o <= x"2000";
when 2308 => read_data_o <= x"2000";
when 2309 => read_data_o <= x"2000";
when 2310 => read_data_o <= x"2000";
when 2311 => read_data_o <= x"2000";
when 2312 => read_data_o <= x"2000";
when 2313 => read_data_o <= x"2000";
when 2314 => read_data_o <= x"2000";
when 2315 => read_data_o <= x"2000";
when 2316 => read_data_o <= x"2000";
when 2317 => read_data_o <= x"2000";
when 2318 => read_data_o <= x"2000";
when 2319 => read_data_o <= x"2000";
when 2320 => read_data_o <= x"2000";
when 2321 => read_data_o <= x"2000";
when 2322 => read_data_o <= x"2000";
when 2323 => read_data_o <= x"2000";
when 2324 => read_data_o <= x"2000";
when 2325 => read_data_o <= x"2000";
when 2326 => read_data_o <= x"2000";
when 2327 => read_data_o <= x"2000";
when 2328 => read_data_o <= x"2000";
when 2329 => read_data_o <= x"2000";
when 2330 => read_data_o <= x"2000";
when 2331 => read_data_o <= x"2000";
when 2332 => read_data_o <= x"2000";
when 2333 => read_data_o <= x"2000";
when 2334 => read_data_o <= x"2000";
when 2335 => read_data_o <= x"2000";
when 2336 => read_data_o <= x"2000";
when 2337 => read_data_o <= x"2000";
when 2338 => read_data_o <= x"2000";
when 2339 => read_data_o <= x"2000";
when 2340 => read_data_o <= x"2000";
when 2341 => read_data_o <= x"2000";
when 2342 => read_data_o <= x"2000";
when 2343 => read_data_o <= x"2000";
when 2344 => read_data_o <= x"2000";
when 2345 => read_data_o <= x"2000";
when 2346 => read_data_o <= x"2000";
when 2347 => read_data_o <= x"2000";
when 2348 => read_data_o <= x"2000";
when 2349 => read_data_o <= x"2000";
when 2350 => read_data_o <= x"2000";
when 2351 => read_data_o <= x"2000";
when 2352 => read_data_o <= x"2000";
when 2353 => read_data_o <= x"2000";
when 2354 => read_data_o <= x"2000";
when 2355 => read_data_o <= x"2000";
when 2356 => read_data_o <= x"2000";
when 2357 => read_data_o <= x"2000";
when 2358 => read_data_o <= x"2000";
when 2359 => read_data_o <= x"2000";
when 2360 => read_data_o <= x"2000";
when 2361 => read_data_o <= x"2000";
when 2362 => read_data_o <= x"2000";
when 2363 => read_data_o <= x"2000";
when 2364 => read_data_o <= x"2000";
when 2365 => read_data_o <= x"2000";
when 2366 => read_data_o <= x"2000";
when 2367 => read_data_o <= x"2000";
when 2368 => read_data_o <= x"2000";
when 2369 => read_data_o <= x"2000";
when 2370 => read_data_o <= x"2000";
when 2371 => read_data_o <= x"2000";
when 2372 => read_data_o <= x"2000";
when 2373 => read_data_o <= x"2000";
when 2374 => read_data_o <= x"2000";
when 2375 => read_data_o <= x"2000";
when 2376 => read_data_o <= x"2000";
when 2377 => read_data_o <= x"2000";
when 2378 => read_data_o <= x"2000";
when 2379 => read_data_o <= x"2000";
when 2380 => read_data_o <= x"2000";
when 2381 => read_data_o <= x"2000";
when 2382 => read_data_o <= x"2000";
when 2383 => read_data_o <= x"2000";
when 2384 => read_data_o <= x"2000";
when 2385 => read_data_o <= x"2000";
when 2386 => read_data_o <= x"2000";
when 2387 => read_data_o <= x"2000";
when 2388 => read_data_o <= x"2000";
when 2389 => read_data_o <= x"2000";
when 2390 => read_data_o <= x"2000";
when 2391 => read_data_o <= x"2000";
when 2392 => read_data_o <= x"2000";
when 2393 => read_data_o <= x"2000";
when 2394 => read_data_o <= x"2000";
when 2395 => read_data_o <= x"2000";
when 2396 => read_data_o <= x"2000";
when 2397 => read_data_o <= x"2000";
when 2398 => read_data_o <= x"2000";
when 2399 => read_data_o <= x"2000";
when 2400 => read_data_o <= x"2000";
when 2401 => read_data_o <= x"2000";
when 2402 => read_data_o <= x"2000";
when 2403 => read_data_o <= x"2000";
when 2404 => read_data_o <= x"2000";
when 2405 => read_data_o <= x"2000";
when 2406 => read_data_o <= x"2000";
when 2407 => read_data_o <= x"2000";
when 2408 => read_data_o <= x"2000";
when 2409 => read_data_o <= x"2000";
when 2410 => read_data_o <= x"2000";
when 2411 => read_data_o <= x"2000";
when 2412 => read_data_o <= x"2000";
when 2413 => read_data_o <= x"2000";
when 2414 => read_data_o <= x"2000";
when 2415 => read_data_o <= x"2000";
when 2416 => read_data_o <= x"2000";
when 2417 => read_data_o <= x"2000";
when 2418 => read_data_o <= x"2000";
when 2419 => read_data_o <= x"2000";
when 2420 => read_data_o <= x"2000";
when 2421 => read_data_o <= x"2000";
when 2422 => read_data_o <= x"2000";
when 2423 => read_data_o <= x"2000";
when 2424 => read_data_o <= x"2000";
when 2425 => read_data_o <= x"2000";
when 2426 => read_data_o <= x"2000";
when 2427 => read_data_o <= x"2000";
when 2428 => read_data_o <= x"2000";
when 2429 => read_data_o <= x"2000";
when 2430 => read_data_o <= x"2000";
when 2431 => read_data_o <= x"2000";
when 2432 => read_data_o <= x"2000";
when 2433 => read_data_o <= x"2000";
when 2434 => read_data_o <= x"2000";
when 2435 => read_data_o <= x"2000";
when 2436 => read_data_o <= x"2000";
when 2437 => read_data_o <= x"2000";
when 2438 => read_data_o <= x"2000";
when 2439 => read_data_o <= x"2000";
when 2440 => read_data_o <= x"2000";
when 2441 => read_data_o <= x"2000";
when 2442 => read_data_o <= x"2000";
when 2443 => read_data_o <= x"2000";
when 2444 => read_data_o <= x"2000";
when 2445 => read_data_o <= x"2000";
when 2446 => read_data_o <= x"2000";
when 2447 => read_data_o <= x"2000";
when 2448 => read_data_o <= x"2000";
when 2449 => read_data_o <= x"2000";
when 2450 => read_data_o <= x"2000";
when 2451 => read_data_o <= x"2000";
when 2452 => read_data_o <= x"2000";
when 2453 => read_data_o <= x"2000";
when 2454 => read_data_o <= x"2000";
when 2455 => read_data_o <= x"2000";
when 2456 => read_data_o <= x"2000";
when 2457 => read_data_o <= x"2000";
when 2458 => read_data_o <= x"2000";
when 2459 => read_data_o <= x"2000";
when 2460 => read_data_o <= x"2000";
when 2461 => read_data_o <= x"2000";
when 2462 => read_data_o <= x"2000";
when 2463 => read_data_o <= x"2000";
when 2464 => read_data_o <= x"2000";
when 2465 => read_data_o <= x"2000";
when 2466 => read_data_o <= x"2000";
when 2467 => read_data_o <= x"2000";
when 2468 => read_data_o <= x"2000";
when 2469 => read_data_o <= x"2000";
when 2470 => read_data_o <= x"2000";
when 2471 => read_data_o <= x"2000";
when 2472 => read_data_o <= x"2000";
when 2473 => read_data_o <= x"2000";
when 2474 => read_data_o <= x"2000";
when 2475 => read_data_o <= x"2000";
when 2476 => read_data_o <= x"2000";
when 2477 => read_data_o <= x"2000";
when 2478 => read_data_o <= x"2000";
when 2479 => read_data_o <= x"2000";
when 2480 => read_data_o <= x"2000";
when 2481 => read_data_o <= x"2000";
when 2482 => read_data_o <= x"2000";
when 2483 => read_data_o <= x"2000";
when 2484 => read_data_o <= x"2000";
when 2485 => read_data_o <= x"2000";
when 2486 => read_data_o <= x"2000";
when 2487 => read_data_o <= x"2000";
when 2488 => read_data_o <= x"2000";
when 2489 => read_data_o <= x"2000";
when 2490 => read_data_o <= x"2000";
when 2491 => read_data_o <= x"2000";
when 2492 => read_data_o <= x"2000";
when 2493 => read_data_o <= x"2000";
when 2494 => read_data_o <= x"2000";
when 2495 => read_data_o <= x"2000";
when 2496 => read_data_o <= x"2000";
when 2497 => read_data_o <= x"2000";
when 2498 => read_data_o <= x"2000";
when 2499 => read_data_o <= x"2000";
when 2500 => read_data_o <= x"2000";
when 2501 => read_data_o <= x"2000";
when 2502 => read_data_o <= x"2000";
when 2503 => read_data_o <= x"2000";
when 2504 => read_data_o <= x"2000";
when 2505 => read_data_o <= x"2000";
when 2506 => read_data_o <= x"2000";
when 2507 => read_data_o <= x"2000";
when 2508 => read_data_o <= x"2000";
when 2509 => read_data_o <= x"2000";
when 2510 => read_data_o <= x"2000";
when 2511 => read_data_o <= x"2000";
when 2512 => read_data_o <= x"2000";
when 2513 => read_data_o <= x"2000";
when 2514 => read_data_o <= x"2000";
when 2515 => read_data_o <= x"2000";
when 2516 => read_data_o <= x"2000";
when 2517 => read_data_o <= x"2000";
when 2518 => read_data_o <= x"2000";
when 2519 => read_data_o <= x"2000";
when 2520 => read_data_o <= x"2000";
when 2521 => read_data_o <= x"2000";
when 2522 => read_data_o <= x"2000";
when 2523 => read_data_o <= x"2000";
when 2524 => read_data_o <= x"2000";
when 2525 => read_data_o <= x"2000";
when 2526 => read_data_o <= x"2000";
when 2527 => read_data_o <= x"2000";
when 2528 => read_data_o <= x"2000";
when 2529 => read_data_o <= x"2000";
when 2530 => read_data_o <= x"2000";
when 2531 => read_data_o <= x"2000";
when 2532 => read_data_o <= x"2000";
when 2533 => read_data_o <= x"2000";
when 2534 => read_data_o <= x"2000";
when 2535 => read_data_o <= x"2000";
when 2536 => read_data_o <= x"2000";
when 2537 => read_data_o <= x"2000";
when 2538 => read_data_o <= x"2000";
when 2539 => read_data_o <= x"2000";
when 2540 => read_data_o <= x"2000";
when 2541 => read_data_o <= x"2000";
when 2542 => read_data_o <= x"2000";
when 2543 => read_data_o <= x"2000";
when 2544 => read_data_o <= x"2000";
when 2545 => read_data_o <= x"2000";
when 2546 => read_data_o <= x"2000";
when 2547 => read_data_o <= x"2000";
when 2548 => read_data_o <= x"2000";
when 2549 => read_data_o <= x"2000";
when 2550 => read_data_o <= x"2000";
when 2551 => read_data_o <= x"2000";
when 2552 => read_data_o <= x"2000";
when 2553 => read_data_o <= x"2000";
when 2554 => read_data_o <= x"2000";
when 2555 => read_data_o <= x"2000";
when 2556 => read_data_o <= x"2000";
when 2557 => read_data_o <= x"2000";
when 2558 => read_data_o <= x"2000";
when 2559 => read_data_o <= x"2000";
when 2560 => read_data_o <= x"2000";
when 2561 => read_data_o <= x"2000";
when 2562 => read_data_o <= x"2000";
when 2563 => read_data_o <= x"2000";
when 2564 => read_data_o <= x"2000";
when 2565 => read_data_o <= x"2000";
when 2566 => read_data_o <= x"2000";
when 2567 => read_data_o <= x"2000";
when 2568 => read_data_o <= x"2000";
when 2569 => read_data_o <= x"2000";
when 2570 => read_data_o <= x"2000";
when 2571 => read_data_o <= x"2000";
when 2572 => read_data_o <= x"2000";
when 2573 => read_data_o <= x"2000";
when 2574 => read_data_o <= x"2000";
when 2575 => read_data_o <= x"2000";
when 2576 => read_data_o <= x"2000";
when 2577 => read_data_o <= x"2000";
when 2578 => read_data_o <= x"2000";
when 2579 => read_data_o <= x"2000";
when 2580 => read_data_o <= x"2000";
when 2581 => read_data_o <= x"2000";
when 2582 => read_data_o <= x"2000";
when 2583 => read_data_o <= x"2000";
when 2584 => read_data_o <= x"2000";
when 2585 => read_data_o <= x"2000";
when 2586 => read_data_o <= x"2000";
when 2587 => read_data_o <= x"2000";
when 2588 => read_data_o <= x"2000";
when 2589 => read_data_o <= x"2000";
when 2590 => read_data_o <= x"2000";
when 2591 => read_data_o <= x"2000";
when 2592 => read_data_o <= x"2000";
when 2593 => read_data_o <= x"2000";
when 2594 => read_data_o <= x"2000";
when 2595 => read_data_o <= x"2000";
when 2596 => read_data_o <= x"2000";
when 2597 => read_data_o <= x"2000";
when 2598 => read_data_o <= x"2000";
when 2599 => read_data_o <= x"2000";
when 2600 => read_data_o <= x"2000";
when 2601 => read_data_o <= x"2000";
when 2602 => read_data_o <= x"2000";
when 2603 => read_data_o <= x"2000";
when 2604 => read_data_o <= x"2000";
when 2605 => read_data_o <= x"2000";
when 2606 => read_data_o <= x"2000";
when 2607 => read_data_o <= x"2000";
when 2608 => read_data_o <= x"2000";
when 2609 => read_data_o <= x"2000";
when 2610 => read_data_o <= x"2000";
when 2611 => read_data_o <= x"2000";
when 2612 => read_data_o <= x"2000";
when 2613 => read_data_o <= x"2000";
when 2614 => read_data_o <= x"2000";
when 2615 => read_data_o <= x"2000";
when 2616 => read_data_o <= x"2000";
when 2617 => read_data_o <= x"2000";
when 2618 => read_data_o <= x"2000";
when 2619 => read_data_o <= x"2000";
when 2620 => read_data_o <= x"2000";
when 2621 => read_data_o <= x"2000";
when 2622 => read_data_o <= x"2000";
when 2623 => read_data_o <= x"2000";
when 2624 => read_data_o <= x"2000";
when 2625 => read_data_o <= x"2000";
when 2626 => read_data_o <= x"2000";
when 2627 => read_data_o <= x"2000";
when 2628 => read_data_o <= x"2000";
when 2629 => read_data_o <= x"2000";
when 2630 => read_data_o <= x"2000";
when 2631 => read_data_o <= x"2000";
when 2632 => read_data_o <= x"2000";
when 2633 => read_data_o <= x"2000";
when 2634 => read_data_o <= x"2000";
when 2635 => read_data_o <= x"2000";
when 2636 => read_data_o <= x"2000";
when 2637 => read_data_o <= x"2000";
when 2638 => read_data_o <= x"2000";
when 2639 => read_data_o <= x"2000";
when 2640 => read_data_o <= x"2000";
when 2641 => read_data_o <= x"2000";
when 2642 => read_data_o <= x"2000";
when 2643 => read_data_o <= x"2000";
when 2644 => read_data_o <= x"2000";
when 2645 => read_data_o <= x"2000";
when 2646 => read_data_o <= x"2000";
when 2647 => read_data_o <= x"2000";
when 2648 => read_data_o <= x"2000";
when 2649 => read_data_o <= x"2000";
when 2650 => read_data_o <= x"2000";
when 2651 => read_data_o <= x"2000";
when 2652 => read_data_o <= x"2000";
when 2653 => read_data_o <= x"2000";
when 2654 => read_data_o <= x"2000";
when 2655 => read_data_o <= x"2000";
when 2656 => read_data_o <= x"2000";
when 2657 => read_data_o <= x"2000";
when 2658 => read_data_o <= x"2000";
when 2659 => read_data_o <= x"2000";
when 2660 => read_data_o <= x"2000";
when 2661 => read_data_o <= x"2000";
when 2662 => read_data_o <= x"2000";
when 2663 => read_data_o <= x"2000";
when 2664 => read_data_o <= x"2000";
when 2665 => read_data_o <= x"2000";
when 2666 => read_data_o <= x"2000";
when 2667 => read_data_o <= x"2000";
when 2668 => read_data_o <= x"2000";
when 2669 => read_data_o <= x"2000";
when 2670 => read_data_o <= x"2000";
when 2671 => read_data_o <= x"2000";
when 2672 => read_data_o <= x"2000";
when 2673 => read_data_o <= x"2000";
when 2674 => read_data_o <= x"2000";
when 2675 => read_data_o <= x"2000";
when 2676 => read_data_o <= x"2000";
when 2677 => read_data_o <= x"2000";
when 2678 => read_data_o <= x"2000";
when 2679 => read_data_o <= x"2000";
when 2680 => read_data_o <= x"2000";
when 2681 => read_data_o <= x"2000";
when 2682 => read_data_o <= x"2000";
when 2683 => read_data_o <= x"2000";
when 2684 => read_data_o <= x"2000";
when 2685 => read_data_o <= x"2000";
when 2686 => read_data_o <= x"2000";
when 2687 => read_data_o <= x"2000";
when 2688 => read_data_o <= x"2000";
when 2689 => read_data_o <= x"2000";
when 2690 => read_data_o <= x"2000";
when 2691 => read_data_o <= x"2000";
when 2692 => read_data_o <= x"2000";
when 2693 => read_data_o <= x"2000";
when 2694 => read_data_o <= x"2000";
when 2695 => read_data_o <= x"2000";
when 2696 => read_data_o <= x"2000";
when 2697 => read_data_o <= x"2000";
when 2698 => read_data_o <= x"2000";
when 2699 => read_data_o <= x"2000";
when 2700 => read_data_o <= x"2000";
when 2701 => read_data_o <= x"2000";
when 2702 => read_data_o <= x"2000";
when 2703 => read_data_o <= x"2000";
when 2704 => read_data_o <= x"2000";
when 2705 => read_data_o <= x"2000";
when 2706 => read_data_o <= x"2000";
when 2707 => read_data_o <= x"2000";
when 2708 => read_data_o <= x"2000";
when 2709 => read_data_o <= x"2000";
when 2710 => read_data_o <= x"2000";
when 2711 => read_data_o <= x"2000";
when 2712 => read_data_o <= x"2000";
when 2713 => read_data_o <= x"2000";
when 2714 => read_data_o <= x"2000";
when 2715 => read_data_o <= x"2000";
when 2716 => read_data_o <= x"2000";
when 2717 => read_data_o <= x"2000";
when 2718 => read_data_o <= x"2000";
when 2719 => read_data_o <= x"2000";
when 2720 => read_data_o <= x"2000";
when 2721 => read_data_o <= x"2000";
when 2722 => read_data_o <= x"2000";
when 2723 => read_data_o <= x"2000";
when 2724 => read_data_o <= x"2000";
when 2725 => read_data_o <= x"2000";
when 2726 => read_data_o <= x"2000";
when 2727 => read_data_o <= x"2000";
when 2728 => read_data_o <= x"2000";
when 2729 => read_data_o <= x"2000";
when 2730 => read_data_o <= x"2000";
when 2731 => read_data_o <= x"2000";
when 2732 => read_data_o <= x"2000";
when 2733 => read_data_o <= x"2000";
when 2734 => read_data_o <= x"2000";
when 2735 => read_data_o <= x"2000";
when 2736 => read_data_o <= x"2000";
when 2737 => read_data_o <= x"2000";
when 2738 => read_data_o <= x"2000";
when 2739 => read_data_o <= x"2000";
when 2740 => read_data_o <= x"2000";
when 2741 => read_data_o <= x"2000";
when 2742 => read_data_o <= x"2000";
when 2743 => read_data_o <= x"2000";
when 2744 => read_data_o <= x"2000";
when 2745 => read_data_o <= x"2000";
when 2746 => read_data_o <= x"2000";
when 2747 => read_data_o <= x"2000";
when 2748 => read_data_o <= x"2000";
when 2749 => read_data_o <= x"2000";
when 2750 => read_data_o <= x"2000";
when 2751 => read_data_o <= x"2000";
when 2752 => read_data_o <= x"2000";
when 2753 => read_data_o <= x"2000";
when 2754 => read_data_o <= x"2000";
when 2755 => read_data_o <= x"2000";
when 2756 => read_data_o <= x"2000";
when 2757 => read_data_o <= x"2000";
when 2758 => read_data_o <= x"2000";
when 2759 => read_data_o <= x"2000";
when 2760 => read_data_o <= x"2000";
when 2761 => read_data_o <= x"2000";
when 2762 => read_data_o <= x"2000";
when 2763 => read_data_o <= x"2000";
when 2764 => read_data_o <= x"2000";
when 2765 => read_data_o <= x"2000";
when 2766 => read_data_o <= x"2000";
when 2767 => read_data_o <= x"2000";
when 2768 => read_data_o <= x"2000";
when 2769 => read_data_o <= x"2000";
when 2770 => read_data_o <= x"2000";
when 2771 => read_data_o <= x"2000";
when 2772 => read_data_o <= x"2000";
when 2773 => read_data_o <= x"2000";
when 2774 => read_data_o <= x"2000";
when 2775 => read_data_o <= x"2000";
when 2776 => read_data_o <= x"2000";
when 2777 => read_data_o <= x"2000";
when 2778 => read_data_o <= x"2000";
when 2779 => read_data_o <= x"2000";
when 2780 => read_data_o <= x"2000";
when 2781 => read_data_o <= x"2000";
when 2782 => read_data_o <= x"2000";
when 2783 => read_data_o <= x"2000";
when 2784 => read_data_o <= x"2000";
when 2785 => read_data_o <= x"2000";
when 2786 => read_data_o <= x"2000";
when 2787 => read_data_o <= x"2000";
when 2788 => read_data_o <= x"2000";
when 2789 => read_data_o <= x"2000";
when 2790 => read_data_o <= x"2000";
when 2791 => read_data_o <= x"2000";
when 2792 => read_data_o <= x"2000";
when 2793 => read_data_o <= x"2000";
when 2794 => read_data_o <= x"2000";
when 2795 => read_data_o <= x"2000";
when 2796 => read_data_o <= x"2000";
when 2797 => read_data_o <= x"2000";
when 2798 => read_data_o <= x"2000";
when 2799 => read_data_o <= x"2000";
when 2800 => read_data_o <= x"2000";
when 2801 => read_data_o <= x"2000";
when 2802 => read_data_o <= x"2000";
when 2803 => read_data_o <= x"2000";
when 2804 => read_data_o <= x"2000";
when 2805 => read_data_o <= x"2000";
when 2806 => read_data_o <= x"2000";
when 2807 => read_data_o <= x"2000";
when 2808 => read_data_o <= x"2000";
when 2809 => read_data_o <= x"2000";
when 2810 => read_data_o <= x"2000";
when 2811 => read_data_o <= x"2000";
when 2812 => read_data_o <= x"2000";
when 2813 => read_data_o <= x"2000";
when 2814 => read_data_o <= x"2000";
when 2815 => read_data_o <= x"2000";
when 2816 => read_data_o <= x"2000";
when 2817 => read_data_o <= x"2000";
when 2818 => read_data_o <= x"2000";
when 2819 => read_data_o <= x"2000";
when 2820 => read_data_o <= x"2000";
when 2821 => read_data_o <= x"2000";
when 2822 => read_data_o <= x"2000";
when 2823 => read_data_o <= x"2000";
when 2824 => read_data_o <= x"2000";
when 2825 => read_data_o <= x"2000";
when 2826 => read_data_o <= x"2000";
when 2827 => read_data_o <= x"2000";
when 2828 => read_data_o <= x"2000";
when 2829 => read_data_o <= x"2000";
when 2830 => read_data_o <= x"2000";
when 2831 => read_data_o <= x"2000";
when 2832 => read_data_o <= x"2000";
when 2833 => read_data_o <= x"2000";
when 2834 => read_data_o <= x"2000";
when 2835 => read_data_o <= x"2000";
when 2836 => read_data_o <= x"2000";
when 2837 => read_data_o <= x"2000";
when 2838 => read_data_o <= x"2000";
when 2839 => read_data_o <= x"2000";
when 2840 => read_data_o <= x"2000";
when 2841 => read_data_o <= x"2000";
when 2842 => read_data_o <= x"2000";
when 2843 => read_data_o <= x"2000";
when 2844 => read_data_o <= x"2000";
when 2845 => read_data_o <= x"2000";
when 2846 => read_data_o <= x"2000";
when 2847 => read_data_o <= x"2000";
when 2848 => read_data_o <= x"2000";
when 2849 => read_data_o <= x"2000";
when 2850 => read_data_o <= x"2000";
when 2851 => read_data_o <= x"2000";
when 2852 => read_data_o <= x"2000";
when 2853 => read_data_o <= x"2000";
when 2854 => read_data_o <= x"2000";
when 2855 => read_data_o <= x"2000";
when 2856 => read_data_o <= x"2000";
when 2857 => read_data_o <= x"2000";
when 2858 => read_data_o <= x"2000";
when 2859 => read_data_o <= x"2000";
when 2860 => read_data_o <= x"2000";
when 2861 => read_data_o <= x"2000";
when 2862 => read_data_o <= x"2000";
when 2863 => read_data_o <= x"2000";
when 2864 => read_data_o <= x"2000";
when 2865 => read_data_o <= x"2000";
when 2866 => read_data_o <= x"2000";
when 2867 => read_data_o <= x"2000";
when 2868 => read_data_o <= x"2000";
when 2869 => read_data_o <= x"2000";
when 2870 => read_data_o <= x"2000";
when 2871 => read_data_o <= x"2000";
when 2872 => read_data_o <= x"2000";
when 2873 => read_data_o <= x"2000";
when 2874 => read_data_o <= x"2000";
when 2875 => read_data_o <= x"2000";
when 2876 => read_data_o <= x"2000";
when 2877 => read_data_o <= x"2000";
when 2878 => read_data_o <= x"2000";
when 2879 => read_data_o <= x"2000";
when 2880 => read_data_o <= x"2000";
when 2881 => read_data_o <= x"2000";
when 2882 => read_data_o <= x"2000";
when 2883 => read_data_o <= x"2000";
when 2884 => read_data_o <= x"2000";
when 2885 => read_data_o <= x"2000";
when 2886 => read_data_o <= x"2000";
when 2887 => read_data_o <= x"2000";
when 2888 => read_data_o <= x"2000";
when 2889 => read_data_o <= x"2000";
when 2890 => read_data_o <= x"2000";
when 2891 => read_data_o <= x"2000";
when 2892 => read_data_o <= x"2000";
when 2893 => read_data_o <= x"2000";
when 2894 => read_data_o <= x"2000";
when 2895 => read_data_o <= x"2000";
when 2896 => read_data_o <= x"2000";
when 2897 => read_data_o <= x"2000";
when 2898 => read_data_o <= x"2000";
when 2899 => read_data_o <= x"2000";
when 2900 => read_data_o <= x"2000";
when 2901 => read_data_o <= x"2000";
when 2902 => read_data_o <= x"2000";
when 2903 => read_data_o <= x"2000";
when 2904 => read_data_o <= x"2000";
when 2905 => read_data_o <= x"2000";
when 2906 => read_data_o <= x"2000";
when 2907 => read_data_o <= x"2000";
when 2908 => read_data_o <= x"2000";
when 2909 => read_data_o <= x"2000";
when 2910 => read_data_o <= x"2000";
when 2911 => read_data_o <= x"2000";
when 2912 => read_data_o <= x"2000";
when 2913 => read_data_o <= x"2000";
when 2914 => read_data_o <= x"2000";
when 2915 => read_data_o <= x"2000";
when 2916 => read_data_o <= x"2000";
when 2917 => read_data_o <= x"2000";
when 2918 => read_data_o <= x"2000";
when 2919 => read_data_o <= x"2000";
when 2920 => read_data_o <= x"2000";
when 2921 => read_data_o <= x"2000";
when 2922 => read_data_o <= x"2000";
when 2923 => read_data_o <= x"2000";
when 2924 => read_data_o <= x"2000";
when 2925 => read_data_o <= x"2000";
when 2926 => read_data_o <= x"2000";
when 2927 => read_data_o <= x"2000";
when 2928 => read_data_o <= x"2000";
when 2929 => read_data_o <= x"2000";
when 2930 => read_data_o <= x"2000";
when 2931 => read_data_o <= x"2000";
when 2932 => read_data_o <= x"2000";
when 2933 => read_data_o <= x"2000";
when 2934 => read_data_o <= x"2000";
when 2935 => read_data_o <= x"2000";
when 2936 => read_data_o <= x"2000";
when 2937 => read_data_o <= x"2000";
when 2938 => read_data_o <= x"2000";
when 2939 => read_data_o <= x"2000";
when 2940 => read_data_o <= x"2000";
when 2941 => read_data_o <= x"2000";
when 2942 => read_data_o <= x"2000";
when 2943 => read_data_o <= x"2000";
when 2944 => read_data_o <= x"2000";
when 2945 => read_data_o <= x"2000";
when 2946 => read_data_o <= x"2000";
when 2947 => read_data_o <= x"2000";
when 2948 => read_data_o <= x"2000";
when 2949 => read_data_o <= x"2000";
when 2950 => read_data_o <= x"2000";
when 2951 => read_data_o <= x"2000";
when 2952 => read_data_o <= x"2000";
when 2953 => read_data_o <= x"2000";
when 2954 => read_data_o <= x"2000";
when 2955 => read_data_o <= x"2000";
when 2956 => read_data_o <= x"2000";
when 2957 => read_data_o <= x"2000";
when 2958 => read_data_o <= x"2000";
when 2959 => read_data_o <= x"2000";
when 2960 => read_data_o <= x"2000";
when 2961 => read_data_o <= x"2000";
when 2962 => read_data_o <= x"2000";
when 2963 => read_data_o <= x"2000";
when 2964 => read_data_o <= x"2000";
when 2965 => read_data_o <= x"2000";
when 2966 => read_data_o <= x"2000";
when 2967 => read_data_o <= x"2000";
when 2968 => read_data_o <= x"2000";
when 2969 => read_data_o <= x"2000";
when 2970 => read_data_o <= x"2000";
when 2971 => read_data_o <= x"2000";
when 2972 => read_data_o <= x"2000";
when 2973 => read_data_o <= x"2000";
when 2974 => read_data_o <= x"2000";
when 2975 => read_data_o <= x"2000";
when 2976 => read_data_o <= x"2000";
when 2977 => read_data_o <= x"2000";
when 2978 => read_data_o <= x"2000";
when 2979 => read_data_o <= x"2000";
when 2980 => read_data_o <= x"2000";
when 2981 => read_data_o <= x"2000";
when 2982 => read_data_o <= x"2000";
when 2983 => read_data_o <= x"2000";
when 2984 => read_data_o <= x"2000";
when 2985 => read_data_o <= x"2000";
when 2986 => read_data_o <= x"2000";
when 2987 => read_data_o <= x"2000";
when 2988 => read_data_o <= x"2000";
when 2989 => read_data_o <= x"2000";
when 2990 => read_data_o <= x"2000";
when 2991 => read_data_o <= x"2000";
when 2992 => read_data_o <= x"2000";
when 2993 => read_data_o <= x"2000";
when 2994 => read_data_o <= x"2000";
when 2995 => read_data_o <= x"2000";
when 2996 => read_data_o <= x"2000";
when 2997 => read_data_o <= x"2000";
when 2998 => read_data_o <= x"2000";
when 2999 => read_data_o <= x"2000";
when 3000 => read_data_o <= x"2000";
when 3001 => read_data_o <= x"2000";
when 3002 => read_data_o <= x"2000";
when 3003 => read_data_o <= x"2000";
when 3004 => read_data_o <= x"2000";
when 3005 => read_data_o <= x"2000";
when 3006 => read_data_o <= x"2000";
when 3007 => read_data_o <= x"2000";
when 3008 => read_data_o <= x"2000";
when 3009 => read_data_o <= x"2000";
when 3010 => read_data_o <= x"2000";
when 3011 => read_data_o <= x"2000";
when 3012 => read_data_o <= x"2000";
when 3013 => read_data_o <= x"2000";
when 3014 => read_data_o <= x"2000";
when 3015 => read_data_o <= x"2000";
when 3016 => read_data_o <= x"2000";
when 3017 => read_data_o <= x"2000";
when 3018 => read_data_o <= x"2000";
when 3019 => read_data_o <= x"2000";
when 3020 => read_data_o <= x"2000";
when 3021 => read_data_o <= x"2000";
when 3022 => read_data_o <= x"2000";
when 3023 => read_data_o <= x"2000";
when 3024 => read_data_o <= x"2000";
when 3025 => read_data_o <= x"2000";
when 3026 => read_data_o <= x"2000";
when 3027 => read_data_o <= x"2000";
when 3028 => read_data_o <= x"2000";
when 3029 => read_data_o <= x"2000";
when 3030 => read_data_o <= x"2000";
when 3031 => read_data_o <= x"2000";
when 3032 => read_data_o <= x"2000";
when 3033 => read_data_o <= x"2000";
when 3034 => read_data_o <= x"2000";
when 3035 => read_data_o <= x"2000";
when 3036 => read_data_o <= x"2000";
when 3037 => read_data_o <= x"2000";
when 3038 => read_data_o <= x"2000";
when 3039 => read_data_o <= x"2000";
when 3040 => read_data_o <= x"2000";
when 3041 => read_data_o <= x"2000";
when 3042 => read_data_o <= x"2000";
when 3043 => read_data_o <= x"2000";
when 3044 => read_data_o <= x"2000";
when 3045 => read_data_o <= x"2000";
when 3046 => read_data_o <= x"2000";
when 3047 => read_data_o <= x"2000";
when 3048 => read_data_o <= x"2000";
when 3049 => read_data_o <= x"2000";
when 3050 => read_data_o <= x"2000";
when 3051 => read_data_o <= x"2000";
when 3052 => read_data_o <= x"2000";
when 3053 => read_data_o <= x"2000";
when 3054 => read_data_o <= x"2000";
when 3055 => read_data_o <= x"2000";
when 3056 => read_data_o <= x"2000";
when 3057 => read_data_o <= x"2000";
when 3058 => read_data_o <= x"2000";
when 3059 => read_data_o <= x"2000";
when 3060 => read_data_o <= x"2000";
when 3061 => read_data_o <= x"2000";
when 3062 => read_data_o <= x"2000";
when 3063 => read_data_o <= x"2000";
when 3064 => read_data_o <= x"2000";
when 3065 => read_data_o <= x"2000";
when 3066 => read_data_o <= x"2000";
when 3067 => read_data_o <= x"2000";
when 3068 => read_data_o <= x"2000";
when 3069 => read_data_o <= x"2000";
when 3070 => read_data_o <= x"2000";
when 3071 => read_data_o <= x"2000";
when 3072 => read_data_o <= x"2000";
when 3073 => read_data_o <= x"2000";
when 3074 => read_data_o <= x"2000";
when 3075 => read_data_o <= x"2000";
when 3076 => read_data_o <= x"2000";
when 3077 => read_data_o <= x"2000";
when 3078 => read_data_o <= x"2000";
when 3079 => read_data_o <= x"2000";
when 3080 => read_data_o <= x"2000";
when 3081 => read_data_o <= x"2000";
when 3082 => read_data_o <= x"2000";
when 3083 => read_data_o <= x"2000";
when 3084 => read_data_o <= x"2000";
when 3085 => read_data_o <= x"2000";
when 3086 => read_data_o <= x"2000";
when 3087 => read_data_o <= x"2000";
when 3088 => read_data_o <= x"2000";
when 3089 => read_data_o <= x"2000";
when 3090 => read_data_o <= x"2000";
when 3091 => read_data_o <= x"2000";
when 3092 => read_data_o <= x"2000";
when 3093 => read_data_o <= x"2000";
when 3094 => read_data_o <= x"2000";
when 3095 => read_data_o <= x"2000";
when 3096 => read_data_o <= x"2000";
when 3097 => read_data_o <= x"2000";
when 3098 => read_data_o <= x"2000";
when 3099 => read_data_o <= x"2000";
when 3100 => read_data_o <= x"2000";
when 3101 => read_data_o <= x"2000";
when 3102 => read_data_o <= x"2000";
when 3103 => read_data_o <= x"2000";
when 3104 => read_data_o <= x"2000";
when 3105 => read_data_o <= x"2000";
when 3106 => read_data_o <= x"2000";
when 3107 => read_data_o <= x"2000";
when 3108 => read_data_o <= x"2000";
when 3109 => read_data_o <= x"2000";
when 3110 => read_data_o <= x"2000";
when 3111 => read_data_o <= x"2000";
when 3112 => read_data_o <= x"2000";
when 3113 => read_data_o <= x"2000";
when 3114 => read_data_o <= x"2000";
when 3115 => read_data_o <= x"2000";
when 3116 => read_data_o <= x"2000";
when 3117 => read_data_o <= x"2000";
when 3118 => read_data_o <= x"2000";
when 3119 => read_data_o <= x"2000";
when 3120 => read_data_o <= x"2000";
when 3121 => read_data_o <= x"2000";
when 3122 => read_data_o <= x"2000";
when 3123 => read_data_o <= x"2000";
when 3124 => read_data_o <= x"2000";
when 3125 => read_data_o <= x"2000";
when 3126 => read_data_o <= x"2000";
when 3127 => read_data_o <= x"2000";
when 3128 => read_data_o <= x"2000";
when 3129 => read_data_o <= x"2000";
when 3130 => read_data_o <= x"2000";
when 3131 => read_data_o <= x"2000";
when 3132 => read_data_o <= x"2000";
when 3133 => read_data_o <= x"2000";
when 3134 => read_data_o <= x"2000";
when 3135 => read_data_o <= x"2000";
when 3136 => read_data_o <= x"2000";
when 3137 => read_data_o <= x"2000";
when 3138 => read_data_o <= x"2000";
when 3139 => read_data_o <= x"2000";
when 3140 => read_data_o <= x"2000";
when 3141 => read_data_o <= x"2000";
when 3142 => read_data_o <= x"2000";
when 3143 => read_data_o <= x"2000";
when 3144 => read_data_o <= x"2000";
when 3145 => read_data_o <= x"2000";
when 3146 => read_data_o <= x"2000";
when 3147 => read_data_o <= x"2000";
when 3148 => read_data_o <= x"2000";
when 3149 => read_data_o <= x"2000";
when 3150 => read_data_o <= x"2000";
when 3151 => read_data_o <= x"2000";
when 3152 => read_data_o <= x"2000";
when 3153 => read_data_o <= x"2000";
when 3154 => read_data_o <= x"2000";
when 3155 => read_data_o <= x"2000";
when 3156 => read_data_o <= x"2000";
when 3157 => read_data_o <= x"2000";
when 3158 => read_data_o <= x"2000";
when 3159 => read_data_o <= x"2000";
when 3160 => read_data_o <= x"2000";
when 3161 => read_data_o <= x"2000";
when 3162 => read_data_o <= x"2000";
when 3163 => read_data_o <= x"2000";
when 3164 => read_data_o <= x"2000";
when 3165 => read_data_o <= x"2000";
when 3166 => read_data_o <= x"2000";
when 3167 => read_data_o <= x"2000";
when 3168 => read_data_o <= x"2000";
when 3169 => read_data_o <= x"2000";
when 3170 => read_data_o <= x"2000";
when 3171 => read_data_o <= x"2000";
when 3172 => read_data_o <= x"2000";
when 3173 => read_data_o <= x"2000";
when 3174 => read_data_o <= x"2000";
when 3175 => read_data_o <= x"2000";
when 3176 => read_data_o <= x"2000";
when 3177 => read_data_o <= x"2000";
when 3178 => read_data_o <= x"2000";
when 3179 => read_data_o <= x"2000";
when 3180 => read_data_o <= x"2000";
when 3181 => read_data_o <= x"2000";
when 3182 => read_data_o <= x"2000";
when 3183 => read_data_o <= x"2000";
when 3184 => read_data_o <= x"2000";
when 3185 => read_data_o <= x"2000";
when 3186 => read_data_o <= x"2000";
when 3187 => read_data_o <= x"2000";
when 3188 => read_data_o <= x"2000";
when 3189 => read_data_o <= x"2000";
when 3190 => read_data_o <= x"2000";
when 3191 => read_data_o <= x"2000";
when 3192 => read_data_o <= x"2000";
when 3193 => read_data_o <= x"2000";
when 3194 => read_data_o <= x"2000";
when 3195 => read_data_o <= x"2000";
when 3196 => read_data_o <= x"2000";
when 3197 => read_data_o <= x"2000";
when 3198 => read_data_o <= x"2000";
when 3199 => read_data_o <= x"2000";
when 3200 => read_data_o <= x"2000";
when 3201 => read_data_o <= x"2000";
when 3202 => read_data_o <= x"2000";
when 3203 => read_data_o <= x"2000";
when 3204 => read_data_o <= x"2000";
when 3205 => read_data_o <= x"2000";
when 3206 => read_data_o <= x"2000";
when 3207 => read_data_o <= x"2000";
when 3208 => read_data_o <= x"2000";
when 3209 => read_data_o <= x"2000";
when 3210 => read_data_o <= x"2000";
when 3211 => read_data_o <= x"2000";
when 3212 => read_data_o <= x"2000";
when 3213 => read_data_o <= x"2000";
when 3214 => read_data_o <= x"2000";
when 3215 => read_data_o <= x"2000";
when 3216 => read_data_o <= x"2000";
when 3217 => read_data_o <= x"2000";
when 3218 => read_data_o <= x"2000";
when 3219 => read_data_o <= x"2000";
when 3220 => read_data_o <= x"2000";
when 3221 => read_data_o <= x"2000";
when 3222 => read_data_o <= x"2000";
when 3223 => read_data_o <= x"2000";
when 3224 => read_data_o <= x"2000";
when 3225 => read_data_o <= x"2000";
when 3226 => read_data_o <= x"2000";
when 3227 => read_data_o <= x"2000";
when 3228 => read_data_o <= x"2000";
when 3229 => read_data_o <= x"2000";
when 3230 => read_data_o <= x"2000";
when 3231 => read_data_o <= x"2000";
when 3232 => read_data_o <= x"2000";
when 3233 => read_data_o <= x"2000";
when 3234 => read_data_o <= x"2000";
when 3235 => read_data_o <= x"2000";
when 3236 => read_data_o <= x"2000";
when 3237 => read_data_o <= x"2000";
when 3238 => read_data_o <= x"2000";
when 3239 => read_data_o <= x"2000";
when 3240 => read_data_o <= x"2000";
when 3241 => read_data_o <= x"2000";
when 3242 => read_data_o <= x"2000";
when 3243 => read_data_o <= x"2000";
when 3244 => read_data_o <= x"2000";
when 3245 => read_data_o <= x"2000";
when 3246 => read_data_o <= x"2000";
when 3247 => read_data_o <= x"2000";
when 3248 => read_data_o <= x"2000";
when 3249 => read_data_o <= x"2000";
when 3250 => read_data_o <= x"2000";
when 3251 => read_data_o <= x"2000";
when 3252 => read_data_o <= x"2000";
when 3253 => read_data_o <= x"2000";
when 3254 => read_data_o <= x"2000";
when 3255 => read_data_o <= x"2000";
when 3256 => read_data_o <= x"2000";
when 3257 => read_data_o <= x"2000";
when 3258 => read_data_o <= x"2000";
when 3259 => read_data_o <= x"2000";
when 3260 => read_data_o <= x"2000";
when 3261 => read_data_o <= x"2000";
when 3262 => read_data_o <= x"2000";
when 3263 => read_data_o <= x"2000";
when 3264 => read_data_o <= x"2000";
when 3265 => read_data_o <= x"2000";
when 3266 => read_data_o <= x"2000";
when 3267 => read_data_o <= x"2000";
when 3268 => read_data_o <= x"2000";
when 3269 => read_data_o <= x"2000";
when 3270 => read_data_o <= x"2000";
when 3271 => read_data_o <= x"2000";
when 3272 => read_data_o <= x"2000";
when 3273 => read_data_o <= x"2000";
when 3274 => read_data_o <= x"2000";
when 3275 => read_data_o <= x"2000";
when 3276 => read_data_o <= x"2000";
when 3277 => read_data_o <= x"2000";
when 3278 => read_data_o <= x"2000";
when 3279 => read_data_o <= x"2000";
when 3280 => read_data_o <= x"2000";
when 3281 => read_data_o <= x"2000";
when 3282 => read_data_o <= x"2000";
when 3283 => read_data_o <= x"2000";
when 3284 => read_data_o <= x"2000";
when 3285 => read_data_o <= x"2000";
when 3286 => read_data_o <= x"2000";
when 3287 => read_data_o <= x"2000";
when 3288 => read_data_o <= x"2000";
when 3289 => read_data_o <= x"2000";
when 3290 => read_data_o <= x"2000";
when 3291 => read_data_o <= x"2000";
when 3292 => read_data_o <= x"2000";
when 3293 => read_data_o <= x"2000";
when 3294 => read_data_o <= x"2000";
when 3295 => read_data_o <= x"2000";
when 3296 => read_data_o <= x"2000";
when 3297 => read_data_o <= x"2000";
when 3298 => read_data_o <= x"2000";
when 3299 => read_data_o <= x"2000";
when 3300 => read_data_o <= x"2000";
when 3301 => read_data_o <= x"2000";
when 3302 => read_data_o <= x"2000";
when 3303 => read_data_o <= x"2000";
when 3304 => read_data_o <= x"2000";
when 3305 => read_data_o <= x"2000";
when 3306 => read_data_o <= x"2000";
when 3307 => read_data_o <= x"2000";
when 3308 => read_data_o <= x"2000";
when 3309 => read_data_o <= x"2000";
when 3310 => read_data_o <= x"2000";
when 3311 => read_data_o <= x"2000";
when 3312 => read_data_o <= x"2000";
when 3313 => read_data_o <= x"2000";
when 3314 => read_data_o <= x"2000";
when 3315 => read_data_o <= x"2000";
when 3316 => read_data_o <= x"2000";
when 3317 => read_data_o <= x"2000";
when 3318 => read_data_o <= x"2000";
when 3319 => read_data_o <= x"2000";
when 3320 => read_data_o <= x"2000";
when 3321 => read_data_o <= x"2000";
when 3322 => read_data_o <= x"2000";
when 3323 => read_data_o <= x"2000";
when 3324 => read_data_o <= x"2000";
when 3325 => read_data_o <= x"2000";
when 3326 => read_data_o <= x"2000";
when 3327 => read_data_o <= x"a000";
when 3328 => read_data_o <= x"0224";
when 3329 => read_data_o <= x"a000";
when 3330 => read_data_o <= x"7040";
when 3331 => read_data_o <= x"00ec";
when 3332 => read_data_o <= x"d02b";
when 3333 => read_data_o <= x"7040";
when 3334 => read_data_o <= x"00cc";
when 3335 => read_data_o <= x"d02b";
when 3336 => read_data_o <= x"7040";
when 3337 => read_data_o <= x"00ac";
when 3338 => read_data_o <= x"d02b";
when 3339 => read_data_o <= x"7040";
when 3340 => read_data_o <= x"008c";
when 3341 => read_data_o <= x"d02b";
when 3342 => read_data_o <= x"a4d0";
when 3343 => read_data_o <= x"a000";
when 3344 => read_data_o <= x"a000";
when 3345 => read_data_o <= x"a000";
when 3346 => read_data_o <= x"a000";
when 3347 => read_data_o <= x"a000";
when 3348 => read_data_o <= x"a000";
when 3349 => read_data_o <= x"a000";
when 3350 => read_data_o <= x"a000";
when 3351 => read_data_o <= x"a000";
when 3352 => read_data_o <= x"a000";
when 3353 => read_data_o <= x"a000";
when 3354 => read_data_o <= x"a000";
when 3355 => read_data_o <= x"a000";
when 3356 => read_data_o <= x"a000";
when 3357 => read_data_o <= x"a000";
when 3358 => read_data_o <= x"a000";
when 3359 => read_data_o <= x"a000";
when 3360 => read_data_o <= x"a000";
when 3361 => read_data_o <= x"a000";
when 3362 => read_data_o <= x"a000";
when 3363 => read_data_o <= x"a000";
when 3364 => read_data_o <= x"a000";
when 3365 => read_data_o <= x"a000";
when 3366 => read_data_o <= x"a000";
when 3367 => read_data_o <= x"a000";
when 3368 => read_data_o <= x"a000";
when 3369 => read_data_o <= x"a000";
when 3370 => read_data_o <= x"a000";
when 3371 => read_data_o <= x"a000";
when 3372 => read_data_o <= x"a000";
when 3373 => read_data_o <= x"a000";
when 3374 => read_data_o <= x"a000";
when 3375 => read_data_o <= x"a000";
when 3376 => read_data_o <= x"a000";
when 3377 => read_data_o <= x"a000";
when 3378 => read_data_o <= x"a000";
when 3379 => read_data_o <= x"a000";
when 3380 => read_data_o <= x"a000";
when 3381 => read_data_o <= x"a000";
when 3382 => read_data_o <= x"a000";
when 3383 => read_data_o <= x"a000";
when 3384 => read_data_o <= x"a000";
when 3385 => read_data_o <= x"a000";
when 3386 => read_data_o <= x"a000";
when 3387 => read_data_o <= x"a000";
when 3388 => read_data_o <= x"a000";
when 3389 => read_data_o <= x"a000";
when 3390 => read_data_o <= x"a000";
when 3391 => read_data_o <= x"a000";
when 3392 => read_data_o <= x"a000";
when 3393 => read_data_o <= x"a000";
when 3394 => read_data_o <= x"a000";
when 3395 => read_data_o <= x"a000";
when 3396 => read_data_o <= x"a000";
when 3397 => read_data_o <= x"a000";
when 3398 => read_data_o <= x"a000";
when 3399 => read_data_o <= x"a000";
when 3400 => read_data_o <= x"a000";
when 3401 => read_data_o <= x"a000";
when 3402 => read_data_o <= x"a000";
when 3403 => read_data_o <= x"a000";
when 3404 => read_data_o <= x"a000";
when 3405 => read_data_o <= x"a000";
when 3406 => read_data_o <= x"a000";
when 3407 => read_data_o <= x"a000";
when 3408 => read_data_o <= x"a000";
when 3409 => read_data_o <= x"a000";
when 3410 => read_data_o <= x"a000";
when 3411 => read_data_o <= x"a000";
when 3412 => read_data_o <= x"a000";
when 3413 => read_data_o <= x"a000";
when 3414 => read_data_o <= x"a000";
when 3415 => read_data_o <= x"a000";
when 3416 => read_data_o <= x"a000";
when 3417 => read_data_o <= x"a000";
when 3418 => read_data_o <= x"a000";
when 3419 => read_data_o <= x"a000";
when 3420 => read_data_o <= x"a000";
when 3421 => read_data_o <= x"a000";
when 3422 => read_data_o <= x"a000";
when 3423 => read_data_o <= x"a000";
when 3424 => read_data_o <= x"a000";
when 3425 => read_data_o <= x"a000";
when 3426 => read_data_o <= x"a000";
when 3427 => read_data_o <= x"a000";
when 3428 => read_data_o <= x"a000";
when 3429 => read_data_o <= x"a000";
when 3430 => read_data_o <= x"a000";
when 3431 => read_data_o <= x"a000";
when 3432 => read_data_o <= x"a000";
when 3433 => read_data_o <= x"a000";
when 3434 => read_data_o <= x"a000";
when 3435 => read_data_o <= x"a000";
when 3436 => read_data_o <= x"a000";
when 3437 => read_data_o <= x"a000";
when 3438 => read_data_o <= x"a000";
when 3439 => read_data_o <= x"a000";
when 3440 => read_data_o <= x"a000";
when 3441 => read_data_o <= x"a000";
when 3442 => read_data_o <= x"a000";
when 3443 => read_data_o <= x"a000";
when 3444 => read_data_o <= x"a000";
when 3445 => read_data_o <= x"a000";
when 3446 => read_data_o <= x"a000";
when 3447 => read_data_o <= x"a000";
when 3448 => read_data_o <= x"a000";
when 3449 => read_data_o <= x"a000";
when 3450 => read_data_o <= x"a000";
when 3451 => read_data_o <= x"a000";
when 3452 => read_data_o <= x"a000";
when 3453 => read_data_o <= x"a000";
when 3454 => read_data_o <= x"a000";
when 3455 => read_data_o <= x"a000";
when 3456 => read_data_o <= x"a000";
when 3457 => read_data_o <= x"a000";
when 3458 => read_data_o <= x"a000";
when 3459 => read_data_o <= x"a000";
when 3460 => read_data_o <= x"a000";
when 3461 => read_data_o <= x"a000";
when 3462 => read_data_o <= x"a000";
when 3463 => read_data_o <= x"a000";
when 3464 => read_data_o <= x"a000";
when 3465 => read_data_o <= x"a000";
when 3466 => read_data_o <= x"a000";
when 3467 => read_data_o <= x"a000";
when 3468 => read_data_o <= x"a000";
when 3469 => read_data_o <= x"a000";
when 3470 => read_data_o <= x"a000";
when 3471 => read_data_o <= x"a000";
when 3472 => read_data_o <= x"a000";
when 3473 => read_data_o <= x"a000";
when 3474 => read_data_o <= x"a000";
when 3475 => read_data_o <= x"a000";
when 3476 => read_data_o <= x"a000";
when 3477 => read_data_o <= x"a000";
when 3478 => read_data_o <= x"a000";
when 3479 => read_data_o <= x"a000";
when 3480 => read_data_o <= x"a000";
when 3481 => read_data_o <= x"a000";
when 3482 => read_data_o <= x"a000";
when 3483 => read_data_o <= x"a000";
when 3484 => read_data_o <= x"a000";
when 3485 => read_data_o <= x"a000";
when 3486 => read_data_o <= x"a000";
when 3487 => read_data_o <= x"a000";
when 3488 => read_data_o <= x"a000";
when 3489 => read_data_o <= x"a000";
when 3490 => read_data_o <= x"a000";
when 3491 => read_data_o <= x"a000";
when 3492 => read_data_o <= x"a000";
when 3493 => read_data_o <= x"a000";
when 3494 => read_data_o <= x"a000";
when 3495 => read_data_o <= x"a000";
when 3496 => read_data_o <= x"a000";
when 3497 => read_data_o <= x"a000";
when 3498 => read_data_o <= x"a000";
when 3499 => read_data_o <= x"a000";
when 3500 => read_data_o <= x"a000";
when 3501 => read_data_o <= x"a000";
when 3502 => read_data_o <= x"a000";
when 3503 => read_data_o <= x"a000";
when 3504 => read_data_o <= x"a000";
when 3505 => read_data_o <= x"a000";
when 3506 => read_data_o <= x"a000";
when 3507 => read_data_o <= x"a000";
when 3508 => read_data_o <= x"a000";
when 3509 => read_data_o <= x"a000";
when 3510 => read_data_o <= x"a000";
when 3511 => read_data_o <= x"a000";
when 3512 => read_data_o <= x"a000";
when 3513 => read_data_o <= x"a000";
when 3514 => read_data_o <= x"a000";
when 3515 => read_data_o <= x"a000";
when 3516 => read_data_o <= x"a000";
when 3517 => read_data_o <= x"a000";
when 3518 => read_data_o <= x"a000";
when 3519 => read_data_o <= x"a000";
when 3520 => read_data_o <= x"a000";
when 3521 => read_data_o <= x"a000";
when 3522 => read_data_o <= x"a000";
when 3523 => read_data_o <= x"a000";
when 3524 => read_data_o <= x"a000";
when 3525 => read_data_o <= x"a000";
when 3526 => read_data_o <= x"a000";
when 3527 => read_data_o <= x"a000";
when 3528 => read_data_o <= x"a000";
when 3529 => read_data_o <= x"a000";
when 3530 => read_data_o <= x"a000";
when 3531 => read_data_o <= x"a000";
when 3532 => read_data_o <= x"a000";
when 3533 => read_data_o <= x"a000";
when 3534 => read_data_o <= x"a000";
when 3535 => read_data_o <= x"a000";
when 3536 => read_data_o <= x"a000";
when 3537 => read_data_o <= x"a000";
when 3538 => read_data_o <= x"a000";
when 3539 => read_data_o <= x"a000";
when 3540 => read_data_o <= x"a000";
when 3541 => read_data_o <= x"a000";
when 3542 => read_data_o <= x"a000";
when 3543 => read_data_o <= x"a000";
when 3544 => read_data_o <= x"a000";
when 3545 => read_data_o <= x"a000";
when 3546 => read_data_o <= x"a000";
when 3547 => read_data_o <= x"a000";
when 3548 => read_data_o <= x"a000";
when 3549 => read_data_o <= x"a000";
when 3550 => read_data_o <= x"a000";
when 3551 => read_data_o <= x"a000";
when 3552 => read_data_o <= x"a000";
when 3553 => read_data_o <= x"a000";
when 3554 => read_data_o <= x"a000";
when 3555 => read_data_o <= x"a000";
when 3556 => read_data_o <= x"a000";
when 3557 => read_data_o <= x"a000";
when 3558 => read_data_o <= x"a000";
when 3559 => read_data_o <= x"a000";
when 3560 => read_data_o <= x"a000";
when 3561 => read_data_o <= x"a000";
when 3562 => read_data_o <= x"a000";
when 3563 => read_data_o <= x"a000";
when 3564 => read_data_o <= x"a000";
when 3565 => read_data_o <= x"a000";
when 3566 => read_data_o <= x"a000";
when 3567 => read_data_o <= x"a000";
when 3568 => read_data_o <= x"a000";
when 3569 => read_data_o <= x"a000";
when 3570 => read_data_o <= x"a000";
when 3571 => read_data_o <= x"a000";
when 3572 => read_data_o <= x"a000";
when 3573 => read_data_o <= x"a000";
when 3574 => read_data_o <= x"a000";
when 3575 => read_data_o <= x"a000";
when 3576 => read_data_o <= x"a000";
when 3577 => read_data_o <= x"a000";
when 3578 => read_data_o <= x"a000";
when 3579 => read_data_o <= x"a000";
when 3580 => read_data_o <= x"a000";
when 3581 => read_data_o <= x"a000";
when 3582 => read_data_o <= x"a000";
when 3583 => read_data_o <= x"a000";
when 3584 => read_data_o <= x"a000";
when 3585 => read_data_o <= x"a000";
when 3586 => read_data_o <= x"a000";
when 3587 => read_data_o <= x"a000";
when 3588 => read_data_o <= x"a000";
when 3589 => read_data_o <= x"a000";
when 3590 => read_data_o <= x"a000";
when 3591 => read_data_o <= x"a000";
when 3592 => read_data_o <= x"a000";
when 3593 => read_data_o <= x"a000";
when 3594 => read_data_o <= x"a000";
when 3595 => read_data_o <= x"a000";
when 3596 => read_data_o <= x"a000";
when 3597 => read_data_o <= x"a000";
when 3598 => read_data_o <= x"a000";
when 3599 => read_data_o <= x"a000";
when 3600 => read_data_o <= x"a000";
when 3601 => read_data_o <= x"a000";
when 3602 => read_data_o <= x"a000";
when 3603 => read_data_o <= x"a000";
when 3604 => read_data_o <= x"a000";
when 3605 => read_data_o <= x"a000";
when 3606 => read_data_o <= x"a000";
when 3607 => read_data_o <= x"a000";
when 3608 => read_data_o <= x"a000";
when 3609 => read_data_o <= x"a000";
when 3610 => read_data_o <= x"a000";
when 3611 => read_data_o <= x"a000";
when 3612 => read_data_o <= x"a000";
when 3613 => read_data_o <= x"a000";
when 3614 => read_data_o <= x"a000";
when 3615 => read_data_o <= x"a000";
when 3616 => read_data_o <= x"a000";
when 3617 => read_data_o <= x"a000";
when 3618 => read_data_o <= x"a000";
when 3619 => read_data_o <= x"a000";
when 3620 => read_data_o <= x"a000";
when 3621 => read_data_o <= x"a000";
when 3622 => read_data_o <= x"a000";
when 3623 => read_data_o <= x"a000";
when 3624 => read_data_o <= x"a000";
when 3625 => read_data_o <= x"a000";
when 3626 => read_data_o <= x"a000";
when 3627 => read_data_o <= x"a000";
when 3628 => read_data_o <= x"a000";
when 3629 => read_data_o <= x"a000";
when 3630 => read_data_o <= x"a000";
when 3631 => read_data_o <= x"a000";
when 3632 => read_data_o <= x"a000";
when 3633 => read_data_o <= x"a000";
when 3634 => read_data_o <= x"a000";
when 3635 => read_data_o <= x"a000";
when 3636 => read_data_o <= x"a000";
when 3637 => read_data_o <= x"a000";
when 3638 => read_data_o <= x"a000";
when 3639 => read_data_o <= x"a000";
when 3640 => read_data_o <= x"a000";
when 3641 => read_data_o <= x"a000";
when 3642 => read_data_o <= x"a000";
when 3643 => read_data_o <= x"a000";
when 3644 => read_data_o <= x"a000";
when 3645 => read_data_o <= x"a000";
when 3646 => read_data_o <= x"a000";
when 3647 => read_data_o <= x"a000";
when 3648 => read_data_o <= x"a000";
when 3649 => read_data_o <= x"a000";
when 3650 => read_data_o <= x"a000";
when 3651 => read_data_o <= x"a000";
when 3652 => read_data_o <= x"a000";
when 3653 => read_data_o <= x"a000";
when 3654 => read_data_o <= x"a000";
when 3655 => read_data_o <= x"a000";
when 3656 => read_data_o <= x"a000";
when 3657 => read_data_o <= x"a000";
when 3658 => read_data_o <= x"a000";
when 3659 => read_data_o <= x"a000";
when 3660 => read_data_o <= x"a000";
when 3661 => read_data_o <= x"a000";
when 3662 => read_data_o <= x"a000";
when 3663 => read_data_o <= x"a000";
when 3664 => read_data_o <= x"a000";
when 3665 => read_data_o <= x"a000";
when 3666 => read_data_o <= x"a000";
when 3667 => read_data_o <= x"a000";
when 3668 => read_data_o <= x"a000";
when 3669 => read_data_o <= x"a000";
when 3670 => read_data_o <= x"a000";
when 3671 => read_data_o <= x"a000";
when 3672 => read_data_o <= x"a000";
when 3673 => read_data_o <= x"a000";
when 3674 => read_data_o <= x"a000";
when 3675 => read_data_o <= x"a000";
when 3676 => read_data_o <= x"a000";
when 3677 => read_data_o <= x"a000";
when 3678 => read_data_o <= x"a000";
when 3679 => read_data_o <= x"a000";
when 3680 => read_data_o <= x"a000";
when 3681 => read_data_o <= x"a000";
when 3682 => read_data_o <= x"a000";
when 3683 => read_data_o <= x"a000";
when 3684 => read_data_o <= x"a000";
when 3685 => read_data_o <= x"a000";
when 3686 => read_data_o <= x"a000";
when 3687 => read_data_o <= x"a000";
when 3688 => read_data_o <= x"a000";
when 3689 => read_data_o <= x"a000";
when 3690 => read_data_o <= x"a000";
when 3691 => read_data_o <= x"a000";
when 3692 => read_data_o <= x"a000";
when 3693 => read_data_o <= x"a000";
when 3694 => read_data_o <= x"a000";
when 3695 => read_data_o <= x"a000";
when 3696 => read_data_o <= x"a000";
when 3697 => read_data_o <= x"a000";
when 3698 => read_data_o <= x"a000";
when 3699 => read_data_o <= x"a000";
when 3700 => read_data_o <= x"a000";
when 3701 => read_data_o <= x"a000";
when 3702 => read_data_o <= x"a000";
when 3703 => read_data_o <= x"a000";
when 3704 => read_data_o <= x"a000";
when 3705 => read_data_o <= x"a000";
when 3706 => read_data_o <= x"a000";
when 3707 => read_data_o <= x"a000";
when 3708 => read_data_o <= x"a000";
when 3709 => read_data_o <= x"a000";
when 3710 => read_data_o <= x"a000";
when 3711 => read_data_o <= x"a000";
when 3712 => read_data_o <= x"a000";
when 3713 => read_data_o <= x"a000";
when 3714 => read_data_o <= x"a000";
when 3715 => read_data_o <= x"a000";
when 3716 => read_data_o <= x"a000";
when 3717 => read_data_o <= x"a000";
when 3718 => read_data_o <= x"a000";
when 3719 => read_data_o <= x"a000";
when 3720 => read_data_o <= x"a000";
when 3721 => read_data_o <= x"a000";
when 3722 => read_data_o <= x"a000";
when 3723 => read_data_o <= x"a000";
when 3724 => read_data_o <= x"a000";
when 3725 => read_data_o <= x"a000";
when 3726 => read_data_o <= x"a000";
when 3727 => read_data_o <= x"a000";
when 3728 => read_data_o <= x"a000";
when 3729 => read_data_o <= x"a000";
when 3730 => read_data_o <= x"a000";
when 3731 => read_data_o <= x"a000";
when 3732 => read_data_o <= x"a000";
when 3733 => read_data_o <= x"a000";
when 3734 => read_data_o <= x"a000";
when 3735 => read_data_o <= x"a000";
when 3736 => read_data_o <= x"a000";
when 3737 => read_data_o <= x"a000";
when 3738 => read_data_o <= x"a000";
when 3739 => read_data_o <= x"a000";
when 3740 => read_data_o <= x"a000";
when 3741 => read_data_o <= x"a000";
when 3742 => read_data_o <= x"a000";
when 3743 => read_data_o <= x"a000";
when 3744 => read_data_o <= x"a000";
when 3745 => read_data_o <= x"a000";
when 3746 => read_data_o <= x"a000";
when 3747 => read_data_o <= x"a000";
when 3748 => read_data_o <= x"a000";
when 3749 => read_data_o <= x"a000";
when 3750 => read_data_o <= x"a000";
when 3751 => read_data_o <= x"a000";
when 3752 => read_data_o <= x"a000";
when 3753 => read_data_o <= x"a000";
when 3754 => read_data_o <= x"a000";
when 3755 => read_data_o <= x"a000";
when 3756 => read_data_o <= x"a000";
when 3757 => read_data_o <= x"a000";
when 3758 => read_data_o <= x"a000";
when 3759 => read_data_o <= x"a000";
when 3760 => read_data_o <= x"a000";
when 3761 => read_data_o <= x"a000";
when 3762 => read_data_o <= x"a000";
when 3763 => read_data_o <= x"a000";
when 3764 => read_data_o <= x"a000";
when 3765 => read_data_o <= x"a000";
when 3766 => read_data_o <= x"a000";
when 3767 => read_data_o <= x"a000";
when 3768 => read_data_o <= x"a000";
when 3769 => read_data_o <= x"a000";
when 3770 => read_data_o <= x"a000";
when 3771 => read_data_o <= x"a000";
when 3772 => read_data_o <= x"a000";
when 3773 => read_data_o <= x"a000";
when 3774 => read_data_o <= x"a000";
when 3775 => read_data_o <= x"a000";
when 3776 => read_data_o <= x"a000";
when 3777 => read_data_o <= x"a000";
when 3778 => read_data_o <= x"a000";
when 3779 => read_data_o <= x"a000";
when 3780 => read_data_o <= x"a000";
when 3781 => read_data_o <= x"a000";
when 3782 => read_data_o <= x"a000";
when 3783 => read_data_o <= x"a000";
when 3784 => read_data_o <= x"a000";
when 3785 => read_data_o <= x"a000";
when 3786 => read_data_o <= x"a000";
when 3787 => read_data_o <= x"a000";
when 3788 => read_data_o <= x"a000";
when 3789 => read_data_o <= x"a000";
when 3790 => read_data_o <= x"a000";
when 3791 => read_data_o <= x"a000";
when 3792 => read_data_o <= x"a000";
when 3793 => read_data_o <= x"a000";
when 3794 => read_data_o <= x"a000";
when 3795 => read_data_o <= x"a000";
when 3796 => read_data_o <= x"a000";
when 3797 => read_data_o <= x"a000";
when 3798 => read_data_o <= x"a000";
when 3799 => read_data_o <= x"a000";
when 3800 => read_data_o <= x"a000";
when 3801 => read_data_o <= x"a000";
when 3802 => read_data_o <= x"a000";
when 3803 => read_data_o <= x"a000";
when 3804 => read_data_o <= x"a000";
when 3805 => read_data_o <= x"a000";
when 3806 => read_data_o <= x"a000";
when 3807 => read_data_o <= x"a000";
when 3808 => read_data_o <= x"a000";
when 3809 => read_data_o <= x"a000";
when 3810 => read_data_o <= x"a000";
when 3811 => read_data_o <= x"a000";
when 3812 => read_data_o <= x"a000";
when 3813 => read_data_o <= x"a000";
when 3814 => read_data_o <= x"a000";
when 3815 => read_data_o <= x"a000";
when 3816 => read_data_o <= x"a000";
when 3817 => read_data_o <= x"a000";
when 3818 => read_data_o <= x"a000";
when 3819 => read_data_o <= x"a000";
when 3820 => read_data_o <= x"a000";
when 3821 => read_data_o <= x"a000";
when 3822 => read_data_o <= x"a000";
when 3823 => read_data_o <= x"a000";
when 3824 => read_data_o <= x"a000";
when 3825 => read_data_o <= x"a000";
when 3826 => read_data_o <= x"a000";
when 3827 => read_data_o <= x"a000";
when 3828 => read_data_o <= x"a000";
when 3829 => read_data_o <= x"a000";
when 3830 => read_data_o <= x"a000";
when 3831 => read_data_o <= x"a000";
when 3832 => read_data_o <= x"a000";
when 3833 => read_data_o <= x"a000";
when 3834 => read_data_o <= x"a000";
when 3835 => read_data_o <= x"a000";
when 3836 => read_data_o <= x"a000";
when 3837 => read_data_o <= x"a000";
when 3838 => read_data_o <= x"a000";
when 3839 => read_data_o <= x"a000";
when 3840 => read_data_o <= x"a000";
when 3841 => read_data_o <= x"a000";
when 3842 => read_data_o <= x"a000";
when 3843 => read_data_o <= x"a000";
when 3844 => read_data_o <= x"a000";
when 3845 => read_data_o <= x"a000";
when 3846 => read_data_o <= x"a000";
when 3847 => read_data_o <= x"a000";
when 3848 => read_data_o <= x"a000";
when 3849 => read_data_o <= x"a000";
when 3850 => read_data_o <= x"a000";
when 3851 => read_data_o <= x"a000";
when 3852 => read_data_o <= x"a000";
when 3853 => read_data_o <= x"a000";
when 3854 => read_data_o <= x"a000";
when 3855 => read_data_o <= x"a000";
when 3856 => read_data_o <= x"a000";
when 3857 => read_data_o <= x"a000";
when 3858 => read_data_o <= x"a000";
when 3859 => read_data_o <= x"a000";
when 3860 => read_data_o <= x"a000";
when 3861 => read_data_o <= x"a000";
when 3862 => read_data_o <= x"a000";
when 3863 => read_data_o <= x"a000";
when 3864 => read_data_o <= x"a000";
when 3865 => read_data_o <= x"a000";
when 3866 => read_data_o <= x"a000";
when 3867 => read_data_o <= x"a000";
when 3868 => read_data_o <= x"a000";
when 3869 => read_data_o <= x"a000";
when 3870 => read_data_o <= x"a000";
when 3871 => read_data_o <= x"a000";
when 3872 => read_data_o <= x"a000";
when 3873 => read_data_o <= x"a000";
when 3874 => read_data_o <= x"a000";
when 3875 => read_data_o <= x"a000";
when 3876 => read_data_o <= x"a000";
when 3877 => read_data_o <= x"a000";
when 3878 => read_data_o <= x"a000";
when 3879 => read_data_o <= x"a000";
when 3880 => read_data_o <= x"a000";
when 3881 => read_data_o <= x"a000";
when 3882 => read_data_o <= x"a000";
when 3883 => read_data_o <= x"a000";
when 3884 => read_data_o <= x"a000";
when 3885 => read_data_o <= x"a000";
when 3886 => read_data_o <= x"a000";
when 3887 => read_data_o <= x"a000";
when 3888 => read_data_o <= x"a000";
when 3889 => read_data_o <= x"a000";
when 3890 => read_data_o <= x"a000";
when 3891 => read_data_o <= x"a000";
when 3892 => read_data_o <= x"a000";
when 3893 => read_data_o <= x"a000";
when 3894 => read_data_o <= x"a000";
when 3895 => read_data_o <= x"a000";
when 3896 => read_data_o <= x"a000";
when 3897 => read_data_o <= x"a000";
when 3898 => read_data_o <= x"a000";
when 3899 => read_data_o <= x"a000";
when 3900 => read_data_o <= x"a000";
when 3901 => read_data_o <= x"a000";
when 3902 => read_data_o <= x"a000";
when 3903 => read_data_o <= x"a000";
when 3904 => read_data_o <= x"a000";
when 3905 => read_data_o <= x"a000";
when 3906 => read_data_o <= x"a000";
when 3907 => read_data_o <= x"a000";
when 3908 => read_data_o <= x"a000";
when 3909 => read_data_o <= x"a000";
when 3910 => read_data_o <= x"a000";
when 3911 => read_data_o <= x"a000";
when 3912 => read_data_o <= x"a000";
when 3913 => read_data_o <= x"a000";
when 3914 => read_data_o <= x"a000";
when 3915 => read_data_o <= x"a000";
when 3916 => read_data_o <= x"a000";
when 3917 => read_data_o <= x"a000";
when 3918 => read_data_o <= x"a000";
when 3919 => read_data_o <= x"a000";
when 3920 => read_data_o <= x"a000";
when 3921 => read_data_o <= x"a000";
when 3922 => read_data_o <= x"a000";
when 3923 => read_data_o <= x"a000";
when 3924 => read_data_o <= x"a000";
when 3925 => read_data_o <= x"a000";
when 3926 => read_data_o <= x"a000";
when 3927 => read_data_o <= x"a000";
when 3928 => read_data_o <= x"a000";
when 3929 => read_data_o <= x"a000";
when 3930 => read_data_o <= x"a000";
when 3931 => read_data_o <= x"a000";
when 3932 => read_data_o <= x"a000";
when 3933 => read_data_o <= x"a000";
when 3934 => read_data_o <= x"a000";
when 3935 => read_data_o <= x"a000";
when 3936 => read_data_o <= x"a000";
when 3937 => read_data_o <= x"a000";
when 3938 => read_data_o <= x"a000";
when 3939 => read_data_o <= x"a000";
when 3940 => read_data_o <= x"a000";
when 3941 => read_data_o <= x"a000";
when 3942 => read_data_o <= x"a000";
when 3943 => read_data_o <= x"a000";
when 3944 => read_data_o <= x"a000";
when 3945 => read_data_o <= x"a000";
when 3946 => read_data_o <= x"a000";
when 3947 => read_data_o <= x"a000";
when 3948 => read_data_o <= x"a000";
when 3949 => read_data_o <= x"a000";
when 3950 => read_data_o <= x"a000";
when 3951 => read_data_o <= x"a000";
when 3952 => read_data_o <= x"a000";
when 3953 => read_data_o <= x"a000";
when 3954 => read_data_o <= x"a000";
when 3955 => read_data_o <= x"a000";
when 3956 => read_data_o <= x"a000";
when 3957 => read_data_o <= x"a000";
when 3958 => read_data_o <= x"a000";
when 3959 => read_data_o <= x"a000";
when 3960 => read_data_o <= x"a000";
when 3961 => read_data_o <= x"a000";
when 3962 => read_data_o <= x"a000";
when 3963 => read_data_o <= x"a000";
when 3964 => read_data_o <= x"a000";
when 3965 => read_data_o <= x"a000";
when 3966 => read_data_o <= x"a000";
when 3967 => read_data_o <= x"a000";
when 3968 => read_data_o <= x"a000";
when 3969 => read_data_o <= x"a000";
when 3970 => read_data_o <= x"a000";
when 3971 => read_data_o <= x"a000";
when 3972 => read_data_o <= x"a000";
when 3973 => read_data_o <= x"a000";
when 3974 => read_data_o <= x"a000";
when 3975 => read_data_o <= x"a000";
when 3976 => read_data_o <= x"a000";
when 3977 => read_data_o <= x"a000";
when 3978 => read_data_o <= x"a000";
when 3979 => read_data_o <= x"a000";
when 3980 => read_data_o <= x"a000";
when 3981 => read_data_o <= x"a000";
when 3982 => read_data_o <= x"a000";
when 3983 => read_data_o <= x"a000";
when 3984 => read_data_o <= x"a000";
when 3985 => read_data_o <= x"a000";
when 3986 => read_data_o <= x"a000";
when 3987 => read_data_o <= x"a000";
when 3988 => read_data_o <= x"a000";
when 3989 => read_data_o <= x"a000";
when 3990 => read_data_o <= x"a000";
when 3991 => read_data_o <= x"a000";
when 3992 => read_data_o <= x"a000";
when 3993 => read_data_o <= x"a000";
when 3994 => read_data_o <= x"a000";
when 3995 => read_data_o <= x"a000";
when 3996 => read_data_o <= x"a000";
when 3997 => read_data_o <= x"a000";
when 3998 => read_data_o <= x"a000";
when 3999 => read_data_o <= x"a000";
when 4000 => read_data_o <= x"a000";
when 4001 => read_data_o <= x"a000";
when 4002 => read_data_o <= x"a000";
when 4003 => read_data_o <= x"a000";
when 4004 => read_data_o <= x"a000";
when 4005 => read_data_o <= x"a000";
when 4006 => read_data_o <= x"a000";
when 4007 => read_data_o <= x"a000";
when 4008 => read_data_o <= x"a000";
when 4009 => read_data_o <= x"a000";
when 4010 => read_data_o <= x"a000";
when 4011 => read_data_o <= x"a000";
when 4012 => read_data_o <= x"a000";
when 4013 => read_data_o <= x"a000";
when 4014 => read_data_o <= x"a000";
when 4015 => read_data_o <= x"a000";
when 4016 => read_data_o <= x"a000";
when 4017 => read_data_o <= x"a000";
when 4018 => read_data_o <= x"a000";
when 4019 => read_data_o <= x"a000";
when 4020 => read_data_o <= x"a000";
when 4021 => read_data_o <= x"a000";
when 4022 => read_data_o <= x"a000";
when 4023 => read_data_o <= x"a000";
when 4024 => read_data_o <= x"a000";
when 4025 => read_data_o <= x"a000";
when 4026 => read_data_o <= x"a000";
when 4027 => read_data_o <= x"a000";
when 4028 => read_data_o <= x"a000";
when 4029 => read_data_o <= x"a000";
when 4030 => read_data_o <= x"a000";
when 4031 => read_data_o <= x"a000";
when 4032 => read_data_o <= x"a000";
when 4033 => read_data_o <= x"a000";
when 4034 => read_data_o <= x"a000";
when 4035 => read_data_o <= x"a000";
when 4036 => read_data_o <= x"a000";
when 4037 => read_data_o <= x"a000";
when 4038 => read_data_o <= x"a000";
when 4039 => read_data_o <= x"a000";
when 4040 => read_data_o <= x"a000";
when 4041 => read_data_o <= x"a000";
when 4042 => read_data_o <= x"a000";
when 4043 => read_data_o <= x"a000";
when 4044 => read_data_o <= x"a000";
when 4045 => read_data_o <= x"a000";
when 4046 => read_data_o <= x"a000";
when 4047 => read_data_o <= x"a000";
when 4048 => read_data_o <= x"a000";
when 4049 => read_data_o <= x"a000";
when 4050 => read_data_o <= x"a000";
when 4051 => read_data_o <= x"a000";
when 4052 => read_data_o <= x"a000";
when 4053 => read_data_o <= x"a000";
when 4054 => read_data_o <= x"a000";
when 4055 => read_data_o <= x"a000";
when 4056 => read_data_o <= x"a000";
when 4057 => read_data_o <= x"a000";
when 4058 => read_data_o <= x"a000";
when 4059 => read_data_o <= x"a000";
when 4060 => read_data_o <= x"a000";
when 4061 => read_data_o <= x"a000";
when 4062 => read_data_o <= x"a000";
when 4063 => read_data_o <= x"a000";
when 4064 => read_data_o <= x"a000";
when 4065 => read_data_o <= x"a000";
when 4066 => read_data_o <= x"a000";
when 4067 => read_data_o <= x"a000";
when 4068 => read_data_o <= x"a000";
when 4069 => read_data_o <= x"a000";
when 4070 => read_data_o <= x"a000";
when 4071 => read_data_o <= x"a000";
when 4072 => read_data_o <= x"a000";
when 4073 => read_data_o <= x"a000";
when 4074 => read_data_o <= x"a000";
when 4075 => read_data_o <= x"a000";
when 4076 => read_data_o <= x"a000";
when 4077 => read_data_o <= x"a000";
when 4078 => read_data_o <= x"a000";
when 4079 => read_data_o <= x"a000";
when 4080 => read_data_o <= x"a000";
when 4081 => read_data_o <= x"a000";
when 4082 => read_data_o <= x"a000";
when 4083 => read_data_o <= x"a000";
when 4084 => read_data_o <= x"a000";
when 4085 => read_data_o <= x"a000";
when 4086 => read_data_o <= x"a000";
when 4087 => read_data_o <= x"a000";
when 4088 => read_data_o <= x"a000";
when 4089 => read_data_o <= x"a000";
when 4090 => read_data_o <= x"a000";
when 4091 => read_data_o <= x"a000";
when 4092 => read_data_o <= x"a000";
when 4093 => read_data_o <= x"a000";
when 4094 => read_data_o <= x"a000";
when 4095 => read_data_o <= x"a000";
when 4096 => read_data_o <= x"6e75";
when 4097 => read_data_o <= x"7665";
when 4098 => read_data_o <= x"6e65";
when 4099 => read_data_o <= x"7473";
when 4100 => read_data_o <= x"44f1";
when 4101 => read_data_o <= x"0000";
when 4102 => read_data_o <= x"0000";
when 4103 => read_data_o <= x"0000";
when 4104 => read_data_o <= x"49e8";
when 4105 => read_data_o <= x"0296";
when 4106 => read_data_o <= x"0000";
when 4107 => read_data_o <= x"0000";
when 4108 => read_data_o <= x"b740";
when 4109 => read_data_o <= x"0353";
when 4110 => read_data_o <= x"0000";
when 4111 => read_data_o <= x"0000";
when 4112 => read_data_o <= x"afa0";
when 4113 => read_data_o <= x"041a";
when 4114 => read_data_o <= x"0000";
when 4115 => read_data_o <= x"0000";
when 4116 => read_data_o <= x"afb0";
when 4117 => read_data_o <= x"041b";
when 4118 => read_data_o <= x"0000";
when 4119 => read_data_o <= x"0000";
when 4120 => read_data_o <= x"0000";
when 4121 => read_data_o <= x"0000";
when 4122 => read_data_o <= x"0000";
when 4123 => read_data_o <= x"0000";
when 4124 => read_data_o <= x"0000";
when 4125 => read_data_o <= x"0000";
when 4126 => read_data_o <= x"0000";
when 4127 => read_data_o <= x"0000";
when 4128 => read_data_o <= x"0000";
when 4129 => read_data_o <= x"0000";
when 4130 => read_data_o <= x"0000";
when 4131 => read_data_o <= x"0000";
when 4132 => read_data_o <= x"d4c8";
when 4133 => read_data_o <= x"041a";
when 4134 => read_data_o <= x"0000";
when 4135 => read_data_o <= x"0000";
when 4136 => read_data_o <= x"0001";
when 4137 => read_data_o <= x"0000";
when 4138 => read_data_o <= x"0000";
when 4139 => read_data_o <= x"0000";
when 4140 => read_data_o <= x"0000";
when 4141 => read_data_o <= x"0000";
when 4142 => read_data_o <= x"0000";
when 4143 => read_data_o <= x"0000";
when 4144 => read_data_o <= x"0000";
when 4145 => read_data_o <= x"0000";
when 4146 => read_data_o <= x"0000";
when 4147 => read_data_o <= x"0000";
when 4148 => read_data_o <= x"0000";
when 4149 => read_data_o <= x"3f80";
when 4150 => read_data_o <= x"6374";
when 4151 => read_data_o <= x"0068";
when 4152 => read_data_o <= x"0000";
when 4153 => read_data_o <= x"0000";
when 4154 => read_data_o <= x"0000";
when 4155 => read_data_o <= x"0000";
when 4156 => read_data_o <= x"0000";
when 4157 => read_data_o <= x"0000";
when 4158 => read_data_o <= x"0000";
when 4159 => read_data_o <= x"0000";
when 4160 => read_data_o <= x"d770";
when 4161 => read_data_o <= x"041a";
when 4162 => read_data_o <= x"0000";
when 4163 => read_data_o <= x"0000";
when 4164 => read_data_o <= x"d770";
when 4165 => read_data_o <= x"041a";
when 4166 => read_data_o <= x"0000";
when 4167 => read_data_o <= x"0000";
when 4168 => read_data_o <= x"0340";
when 4169 => read_data_o <= x"041b";
when 4170 => read_data_o <= x"0000";
when 4171 => read_data_o <= x"0000";
when 4172 => read_data_o <= x"03a8";
when 4173 => read_data_o <= x"041b";
when 4174 => read_data_o <= x"0000";
when 4175 => read_data_o <= x"0000";
when 4176 => read_data_o <= x"2400";
when 4177 => read_data_o <= x"00f4";
when 4178 => read_data_o <= x"2400";
when 4179 => read_data_o <= x"00f4";
when 4180 => read_data_o <= x"2400";
when 4181 => read_data_o <= x"00f4";
when 4182 => read_data_o <= x"0000";
when 4183 => read_data_o <= x"0000";
when 4184 => read_data_o <= x"0000";
when 4185 => read_data_o <= x"0000";
when 4186 => read_data_o <= x"0000";
when 4187 => read_data_o <= x"3ff0";
when 4188 => read_data_o <= x"5100";
when 4189 => read_data_o <= x"8d4a";
when 4190 => read_data_o <= x"000e";
when 4191 => read_data_o <= x"0000";
when 4192 => read_data_o <= x"0000";
when 4193 => read_data_o <= x"0000";
when 4194 => read_data_o <= x"0000";
when 4195 => read_data_o <= x"0000";
when 4196 => read_data_o <= x"ad00";
when 4197 => read_data_o <= x"4d2d";
when 4198 => read_data_o <= x"7fff";
when 4199 => read_data_o <= x"0000";
when 4200 => read_data_o <= x"0000";
when 4201 => read_data_o <= x"0000";
when 4202 => read_data_o <= x"0000";
when 4203 => read_data_o <= x"0000";
when 4204 => read_data_o <= x"0000";
when 4205 => read_data_o <= x"0000";
when 4206 => read_data_o <= x"0000";
when 4207 => read_data_o <= x"0000";
when 4208 => read_data_o <= x"d540";
when 4209 => read_data_o <= x"041a";
when 4210 => read_data_o <= x"0000";
when 4211 => read_data_o <= x"0000";
when 4212 => read_data_o <= x"0000";
when 4213 => read_data_o <= x"0000";
when 4214 => read_data_o <= x"0000";
when 4215 => read_data_o <= x"0000";
when 4216 => read_data_o <= x"0000";
when 4217 => read_data_o <= x"0000";
when 4218 => read_data_o <= x"0000";
when 4219 => read_data_o <= x"0000";
when 4220 => read_data_o <= x"0000";
when 4221 => read_data_o <= x"0000";
when 4222 => read_data_o <= x"0000";
when 4223 => read_data_o <= x"0000";
when 4224 => read_data_o <= x"adb0";
when 4225 => read_data_o <= x"4d2d";
when 4226 => read_data_o <= x"7fff";
when 4227 => read_data_o <= x"0000";
when 4228 => read_data_o <= x"afe0";
when 4229 => read_data_o <= x"4d2d";
when 4230 => read_data_o <= x"7fff";
when 4231 => read_data_o <= x"0000";
when 4232 => read_data_o <= x"d570";
when 4233 => read_data_o <= x"041a";
when 4234 => read_data_o <= x"0000";
when 4235 => read_data_o <= x"0000";
when 4236 => read_data_o <= x"0008";
when 4237 => read_data_o <= x"0000";
when 4238 => read_data_o <= x"0000";
when 4239 => read_data_o <= x"0000";
when 4240 => read_data_o <= x"6d3a";
when 4241 => read_data_o <= x"6961";
when 4242 => read_data_o <= x"636e";
when 4243 => read_data_o <= x"7570";
when 4244 => read_data_o <= x"0000";
when 4245 => read_data_o <= x"0000";
when 4246 => read_data_o <= x"0000";
when 4247 => read_data_o <= x"0000";
when 4248 => read_data_o <= x"d590";
when 4249 => read_data_o <= x"041a";
when 4250 => read_data_o <= x"0000";
when 4251 => read_data_o <= x"0000";
when 4252 => read_data_o <= x"0007";
when 4253 => read_data_o <= x"0000";
when 4254 => read_data_o <= x"0000";
when 4255 => read_data_o <= x"0000";
when 4256 => read_data_o <= x"616d";
when 4257 => read_data_o <= x"6e69";
when 4258 => read_data_o <= x"7063";
when 4259 => read_data_o <= x"0075";
when 4260 => read_data_o <= x"0000";
when 4261 => read_data_o <= x"0000";
when 4262 => read_data_o <= x"0000";
when 4263 => read_data_o <= x"0000";
when 4264 => read_data_o <= x"0101";
when 4265 => read_data_o <= x"0030";
when 4266 => read_data_o <= x"7f00";
when 4267 => read_data_o <= x"0000";
when 4268 => read_data_o <= x"0000";
when 4269 => read_data_o <= x"0000";
when 4270 => read_data_o <= x"0000";
when 4271 => read_data_o <= x"0000";
when 4272 => read_data_o <= x"6ea0";
when 4273 => read_data_o <= x"04be";
when 4274 => read_data_o <= x"0000";
when 4275 => read_data_o <= x"0000";
when 4276 => read_data_o <= x"6ef0";
when 4277 => read_data_o <= x"04be";
when 4278 => read_data_o <= x"0000";
when 4279 => read_data_o <= x"0000";
when 4280 => read_data_o <= x"6ef0";
when 4281 => read_data_o <= x"04be";
when 4282 => read_data_o <= x"0000";
when 4283 => read_data_o <= x"0000";
when 4284 => read_data_o <= x"d5c8";
when 4285 => read_data_o <= x"041a";
when 4286 => read_data_o <= x"0000";
when 4287 => read_data_o <= x"0000";
when 4288 => read_data_o <= x"d5c8";
when 4289 => read_data_o <= x"041a";
when 4290 => read_data_o <= x"0000";
when 4291 => read_data_o <= x"0000";
when 4292 => read_data_o <= x"0000";
when 4293 => read_data_o <= x"0000";
when 4294 => read_data_o <= x"0000";
when 4295 => read_data_o <= x"0000";
when 4296 => read_data_o <= x"0000";
when 4297 => read_data_o <= x"0000";
when 4298 => read_data_o <= x"0000";
when 4299 => read_data_o <= x"0000";
when 4300 => read_data_o <= x"0000";
when 4301 => read_data_o <= x"0000";
when 4302 => read_data_o <= x"0000";
when 4303 => read_data_o <= x"0000";
when 4304 => read_data_o <= x"0000";
when 4305 => read_data_o <= x"0000";
when 4306 => read_data_o <= x"0000";
when 4307 => read_data_o <= x"0000";
when 4308 => read_data_o <= x"f5d8";
when 4309 => read_data_o <= x"02ad";
when 4310 => read_data_o <= x"0000";
when 4311 => read_data_o <= x"0000";
when 4312 => read_data_o <= x"f9c0";
when 4313 => read_data_o <= x"0289";
when 4314 => read_data_o <= x"0000";
when 4315 => read_data_o <= x"0000";
when 4316 => read_data_o <= x"0000";
when 4317 => read_data_o <= x"0000";
when 4318 => read_data_o <= x"0000";
when 4319 => read_data_o <= x"0000";
when 4320 => read_data_o <= x"0000";
when 4321 => read_data_o <= x"0000";
when 4322 => read_data_o <= x"0000";
when 4323 => read_data_o <= x"0000";
when 4324 => read_data_o <= x"0000";
when 4325 => read_data_o <= x"0000";
when 4326 => read_data_o <= x"0000";
when 4327 => read_data_o <= x"0000";
when 4328 => read_data_o <= x"4720";
when 4329 => read_data_o <= x"04b3";
when 4330 => read_data_o <= x"0000";
when 4331 => read_data_o <= x"0000";
when 4332 => read_data_o <= x"4720";
when 4333 => read_data_o <= x"04b3";
when 4334 => read_data_o <= x"0000";
when 4335 => read_data_o <= x"0000";
when 4336 => read_data_o <= x"4b20";
when 4337 => read_data_o <= x"04b3";
when 4338 => read_data_o <= x"0000";
when 4339 => read_data_o <= x"0000";
when 4340 => read_data_o <= x"ed60";
when 4341 => read_data_o <= x"858b";
when 4342 => read_data_o <= x"7f4f";
when 4343 => read_data_o <= x"0000";
when 4344 => read_data_o <= x"0010";
when 4345 => read_data_o <= x"0000";
when 4346 => read_data_o <= x"0000";
when 4347 => read_data_o <= x"0000";
when 4348 => read_data_o <= x"4720";
when 4349 => read_data_o <= x"04b3";
when 4350 => read_data_o <= x"0000";
when 4351 => read_data_o <= x"0000";
when 4352 => read_data_o <= x"4b20";
when 4353 => read_data_o <= x"04b3";
when 4354 => read_data_o <= x"0000";
when 4355 => read_data_o <= x"0000";
when 4356 => read_data_o <= x"4b20";
when 4357 => read_data_o <= x"04b3";
when 4358 => read_data_o <= x"0000";
when 4359 => read_data_o <= x"0000";
when 4360 => read_data_o <= x"4720";
when 4361 => read_data_o <= x"04b3";
when 4362 => read_data_o <= x"0000";
when 4363 => read_data_o <= x"0000";
when 4364 => read_data_o <= x"f600";
when 4365 => read_data_o <= x"02ad";
when 4366 => read_data_o <= x"0000";
when 4367 => read_data_o <= x"0000";
when 4368 => read_data_o <= x"0006";
when 4369 => read_data_o <= x"0000";
when 4370 => read_data_o <= x"0000";
when 4371 => read_data_o <= x"0000";
when 4372 => read_data_o <= x"0000";
when 4373 => read_data_o <= x"0000";
when 4374 => read_data_o <= x"0000";
when 4375 => read_data_o <= x"0000";
when 4376 => read_data_o <= x"1002";
when 4377 => read_data_o <= x"0000";
when 4378 => read_data_o <= x"0000";
when 4379 => read_data_o <= x"0000";
when 4380 => read_data_o <= x"0000";
when 4381 => read_data_o <= x"0000";
when 4382 => read_data_o <= x"0000";
when 4383 => read_data_o <= x"0000";
when 4384 => read_data_o <= x"0000";
when 4385 => read_data_o <= x"0000";
when 4386 => read_data_o <= x"0000";
when 4387 => read_data_o <= x"0000";
when 4388 => read_data_o <= x"0000";
when 4389 => read_data_o <= x"0000";
when 4390 => read_data_o <= x"0000";
when 4391 => read_data_o <= x"0000";
when 4392 => read_data_o <= x"0000";
when 4393 => read_data_o <= x"0000";
when 4394 => read_data_o <= x"0000";
when 4395 => read_data_o <= x"0000";
when 4396 => read_data_o <= x"0000";
when 4397 => read_data_o <= x"0000";
when 4398 => read_data_o <= x"0000";
when 4399 => read_data_o <= x"0000";
when 4400 => read_data_o <= x"0000";
when 4401 => read_data_o <= x"0000";
when 4402 => read_data_o <= x"0000";
when 4403 => read_data_o <= x"0000";
when 4404 => read_data_o <= x"0000";
when 4405 => read_data_o <= x"0000";
when 4406 => read_data_o <= x"0000";
when 4407 => read_data_o <= x"0000";
when 4408 => read_data_o <= x"0000";
when 4409 => read_data_o <= x"0000";
when 4410 => read_data_o <= x"0000";
when 4411 => read_data_o <= x"0000";
when 4412 => read_data_o <= x"0000";
when 4413 => read_data_o <= x"0000";
when 4414 => read_data_o <= x"0000";
when 4415 => read_data_o <= x"0000";
when 4416 => read_data_o <= x"0000";
when 4417 => read_data_o <= x"0000";
when 4418 => read_data_o <= x"0000";
when 4419 => read_data_o <= x"0000";
when 4420 => read_data_o <= x"0000";
when 4421 => read_data_o <= x"0000";
when 4422 => read_data_o <= x"0000";
when 4423 => read_data_o <= x"0000";
when 4424 => read_data_o <= x"0000";
when 4425 => read_data_o <= x"0000";
when 4426 => read_data_o <= x"0000";
when 4427 => read_data_o <= x"0000";
when 4428 => read_data_o <= x"0000";
when 4429 => read_data_o <= x"0000";
when 4430 => read_data_o <= x"0000";
when 4431 => read_data_o <= x"0000";
when 4432 => read_data_o <= x"0000";
when 4433 => read_data_o <= x"0000";
when 4434 => read_data_o <= x"0000";
when 4435 => read_data_o <= x"0000";
when 4436 => read_data_o <= x"0000";
when 4437 => read_data_o <= x"0000";
when 4438 => read_data_o <= x"0000";
when 4439 => read_data_o <= x"0000";
when 4440 => read_data_o <= x"0000";
when 4441 => read_data_o <= x"0000";
when 4442 => read_data_o <= x"0000";
when 4443 => read_data_o <= x"0000";
when 4444 => read_data_o <= x"0000";
when 4445 => read_data_o <= x"0000";
when 4446 => read_data_o <= x"0000";
when 4447 => read_data_o <= x"0000";
when 4448 => read_data_o <= x"0000";
when 4449 => read_data_o <= x"0000";
when 4450 => read_data_o <= x"0000";
when 4451 => read_data_o <= x"0000";
when 4452 => read_data_o <= x"0000";
when 4453 => read_data_o <= x"0000";
when 4454 => read_data_o <= x"0000";
when 4455 => read_data_o <= x"0000";
when 4456 => read_data_o <= x"0000";
when 4457 => read_data_o <= x"0000";
when 4458 => read_data_o <= x"0000";
when 4459 => read_data_o <= x"0000";
when 4460 => read_data_o <= x"0008";
when 4461 => read_data_o <= x"0000";
when 4462 => read_data_o <= x"7968";
when 4463 => read_data_o <= x"0000";
when 4464 => read_data_o <= x"d6a8";
when 4465 => read_data_o <= x"041a";
when 4466 => read_data_o <= x"0000";
when 4467 => read_data_o <= x"0000";
when 4468 => read_data_o <= x"ed60";
when 4469 => read_data_o <= x"858b";
when 4470 => read_data_o <= x"7f4f";
when 4471 => read_data_o <= x"0000";
when 4472 => read_data_o <= x"0000";
when 4473 => read_data_o <= x"0000";
when 4474 => read_data_o <= x"0000";
when 4475 => read_data_o <= x"0000";
when 4476 => read_data_o <= x"0000";
when 4477 => read_data_o <= x"0000";
when 4478 => read_data_o <= x"0000";
when 4479 => read_data_o <= x"0000";
when 4480 => read_data_o <= x"d600";
when 4481 => read_data_o <= x"041a";
when 4482 => read_data_o <= x"0000";
when 4483 => read_data_o <= x"0000";
when 4484 => read_data_o <= x"e780";
when 4485 => read_data_o <= x"858b";
when 4486 => read_data_o <= x"7f4f";
when 4487 => read_data_o <= x"0000";
when 4488 => read_data_o <= x"e710";
when 4489 => read_data_o <= x"858b";
when 4490 => read_data_o <= x"7f4f";
when 4491 => read_data_o <= x"0000";
when 4492 => read_data_o <= x"e720";
when 4493 => read_data_o <= x"858b";
when 4494 => read_data_o <= x"7f4f";
when 4495 => read_data_o <= x"0000";
when 4496 => read_data_o <= x"4af0";
when 4497 => read_data_o <= x"0296";
when 4498 => read_data_o <= x"0000";
when 4499 => read_data_o <= x"0000";
when 4500 => read_data_o <= x"0340";
when 4501 => read_data_o <= x"041b";
when 4502 => read_data_o <= x"0000";
when 4503 => read_data_o <= x"0000";
when 4504 => read_data_o <= x"d460";
when 4505 => read_data_o <= x"041a";
when 4506 => read_data_o <= x"0000";
when 4507 => read_data_o <= x"0000";
when 4508 => read_data_o <= x"5b0a";
when 4509 => read_data_o <= x"0299";
when 4510 => read_data_o <= x"0000";
when 4511 => read_data_o <= x"0000";
when 4512 => read_data_o <= x"0258";
when 4513 => read_data_o <= x"4d2e";
when 4514 => read_data_o <= x"7fff";
when 4515 => read_data_o <= x"0000";
when 4516 => read_data_o <= x"0000";
when 4517 => read_data_o <= x"0000";
when 4518 => read_data_o <= x"0000";
when 4519 => read_data_o <= x"0000";
when 4520 => read_data_o <= x"0000";
when 4521 => read_data_o <= x"0000";
when 4522 => read_data_o <= x"0000";
when 4523 => read_data_o <= x"0000";
when 4524 => read_data_o <= x"0000";
when 4525 => read_data_o <= x"0000";
when 4526 => read_data_o <= x"0000";
when 4527 => read_data_o <= x"0000";
when 4528 => read_data_o <= x"0000";
when 4529 => read_data_o <= x"0000";
when 4530 => read_data_o <= x"0000";
when 4531 => read_data_o <= x"0000";
when 4532 => read_data_o <= x"0000";
when 4533 => read_data_o <= x"0000";
when 4534 => read_data_o <= x"0000";
when 4535 => read_data_o <= x"0000";
when 4536 => read_data_o <= x"0000";
when 4537 => read_data_o <= x"0000";
when 4538 => read_data_o <= x"0000";
when 4539 => read_data_o <= x"0000";
when 4540 => read_data_o <= x"0000";
when 4541 => read_data_o <= x"0000";
when 4542 => read_data_o <= x"0000";
when 4543 => read_data_o <= x"0000";
when 4544 => read_data_o <= x"0000";
when 4545 => read_data_o <= x"0000";
when 4546 => read_data_o <= x"0003";
when 4547 => read_data_o <= x"0000";
when 4548 => read_data_o <= x"2540";
when 4549 => read_data_o <= x"02a7";
when 4550 => read_data_o <= x"0000";
when 4551 => read_data_o <= x"0000";
when 4552 => read_data_o <= x"0000";
when 4553 => read_data_o <= x"0000";
when 4554 => read_data_o <= x"0000";
when 4555 => read_data_o <= x"0000";
when 4556 => read_data_o <= x"0000";
when 4557 => read_data_o <= x"0000";
when 4558 => read_data_o <= x"0000";
when 4559 => read_data_o <= x"0000";
when 4560 => read_data_o <= x"0000";
when 4561 => read_data_o <= x"0000";
when 4562 => read_data_o <= x"0000";
when 4563 => read_data_o <= x"0000";
when 4564 => read_data_o <= x"d460";
when 4565 => read_data_o <= x"041a";
when 4566 => read_data_o <= x"0000";
when 4567 => read_data_o <= x"0000";
when 4568 => read_data_o <= x"0000";
when 4569 => read_data_o <= x"0000";
when 4570 => read_data_o <= x"0000";
when 4571 => read_data_o <= x"0000";
when 4572 => read_data_o <= x"0000";
when 4573 => read_data_o <= x"0000";
when 4574 => read_data_o <= x"0000";
when 4575 => read_data_o <= x"0000";
when 4576 => read_data_o <= x"0000";
when 4577 => read_data_o <= x"0000";
when 4578 => read_data_o <= x"0000";
when 4579 => read_data_o <= x"0000";
when 4580 => read_data_o <= x"0000";
when 4581 => read_data_o <= x"0000";
when 4582 => read_data_o <= x"0000";
when 4583 => read_data_o <= x"0000";
when 4584 => read_data_o <= x"0000";
when 4585 => read_data_o <= x"0000";
when 4586 => read_data_o <= x"0000";
when 4587 => read_data_o <= x"0000";
when 4588 => read_data_o <= x"0000";
when 4589 => read_data_o <= x"0000";
when 4590 => read_data_o <= x"0000";
when 4591 => read_data_o <= x"0000";
when 4592 => read_data_o <= x"0000";
when 4593 => read_data_o <= x"0000";
when 4594 => read_data_o <= x"0000";
when 4595 => read_data_o <= x"0000";
when 4596 => read_data_o <= x"0000";
when 4597 => read_data_o <= x"0000";
when 4598 => read_data_o <= x"6374";
when 4599 => read_data_o <= x"0068";
when 4600 => read_data_o <= x"d850";
when 4601 => read_data_o <= x"041a";
when 4602 => read_data_o <= x"0000";
when 4603 => read_data_o <= x"0000";
when 4604 => read_data_o <= x"0000";
when 4605 => read_data_o <= x"0000";
when 4606 => read_data_o <= x"0000";
when 4607 => read_data_o <= x"0000";
when 4608 => read_data_o <= x"0000";
when 4609 => read_data_o <= x"0000";
when 4610 => read_data_o <= x"0000";
when 4611 => read_data_o <= x"0000";
when 4612 => read_data_o <= x"ff20";
when 4613 => read_data_o <= x"ffff";
when 4614 => read_data_o <= x"ffff";
when 4615 => read_data_o <= x"ffff";
when 4616 => read_data_o <= x"0000";
when 4617 => read_data_o <= x"0000";
when 4618 => read_data_o <= x"0000";
when 4619 => read_data_o <= x"0000";
when 4620 => read_data_o <= x"d460";
when 4621 => read_data_o <= x"041a";
when 4622 => read_data_o <= x"0000";
when 4623 => read_data_o <= x"0000";
when 4624 => read_data_o <= x"0000";
when 4625 => read_data_o <= x"0000";
when 4626 => read_data_o <= x"0000";
when 4627 => read_data_o <= x"0000";
when 4628 => read_data_o <= x"0000";
when 4629 => read_data_o <= x"0000";
when 4630 => read_data_o <= x"7fff";
when 4631 => read_data_o <= x"0000";
when 4632 => read_data_o <= x"0000";
when 4633 => read_data_o <= x"0000";
when 4634 => read_data_o <= x"0000";
when 4635 => read_data_o <= x"0000";
when 4636 => read_data_o <= x"0000";
when 4637 => read_data_o <= x"0000";
when 4638 => read_data_o <= x"0000";
when 4639 => read_data_o <= x"0000";
when 4640 => read_data_o <= x"0000";
when 4641 => read_data_o <= x"0000";
when 4642 => read_data_o <= x"0000";
when 4643 => read_data_o <= x"0000";
when 4644 => read_data_o <= x"0000";
when 4645 => read_data_o <= x"0000";
when 4646 => read_data_o <= x"0000";
when 4647 => read_data_o <= x"0000";
when 4648 => read_data_o <= x"0000";
when 4649 => read_data_o <= x"0000";
when 4650 => read_data_o <= x"0000";
when 4651 => read_data_o <= x"0000";
when 4652 => read_data_o <= x"0000";
when 4653 => read_data_o <= x"0000";
when 4654 => read_data_o <= x"0000";
when 4655 => read_data_o <= x"0000";
when 4656 => read_data_o <= x"0000";
when 4657 => read_data_o <= x"0000";
when 4658 => read_data_o <= x"0000";
when 4659 => read_data_o <= x"0000";
when 4660 => read_data_o <= x"0000";
when 4661 => read_data_o <= x"0000";
when 4662 => read_data_o <= x"d278";
when 4663 => read_data_o <= x"f831";
when 4664 => read_data_o <= x"0000";
when 4665 => read_data_o <= x"0000";
when 4666 => read_data_o <= x"0000";
when 4667 => read_data_o <= x"0000";
when 4668 => read_data_o <= x"0041";
when 4669 => read_data_o <= x"0000";
when 4670 => read_data_o <= x"0000";
when 4671 => read_data_o <= x"0000";
when 4672 => read_data_o <= x"0000";
when 4673 => read_data_o <= x"0000";
when 4674 => read_data_o <= x"0000";
when 4675 => read_data_o <= x"0000";
when 4676 => read_data_o <= x"af90";
when 4677 => read_data_o <= x"041a";
when 4678 => read_data_o <= x"0000";
when 4679 => read_data_o <= x"0000";
when 4680 => read_data_o <= x"0000";
when 4681 => read_data_o <= x"0000";
when 4682 => read_data_o <= x"0000";
when 4683 => read_data_o <= x"0000";
when 4684 => read_data_o <= x"d460";
when 4685 => read_data_o <= x"041a";
when 4686 => read_data_o <= x"0000";
when 4687 => read_data_o <= x"0000";
when 4688 => read_data_o <= x"0000";
when 4689 => read_data_o <= x"0000";
when 4690 => read_data_o <= x"0000";
when 4691 => read_data_o <= x"0000";
when 4692 => read_data_o <= x"d770";
when 4693 => read_data_o <= x"041a";
when 4694 => read_data_o <= x"0000";
when 4695 => read_data_o <= x"0000";
when 4696 => read_data_o <= x"0000";
when 4697 => read_data_o <= x"0000";
when 4698 => read_data_o <= x"0000";
when 4699 => read_data_o <= x"0000";
when 4700 => read_data_o <= x"0000";
when 4701 => read_data_o <= x"0000";
when 4702 => read_data_o <= x"0000";
when 4703 => read_data_o <= x"0000";
when 4704 => read_data_o <= x"0000";
when 4705 => read_data_o <= x"0000";
when 4706 => read_data_o <= x"0000";
when 4707 => read_data_o <= x"0000";
when 4708 => read_data_o <= x"0000";
when 4709 => read_data_o <= x"0000";
when 4710 => read_data_o <= x"0000";
when 4711 => read_data_o <= x"0000";
when 4712 => read_data_o <= x"0000";
when 4713 => read_data_o <= x"0000";
when 4714 => read_data_o <= x"0000";
when 4715 => read_data_o <= x"0000";
when 4716 => read_data_o <= x"0000";
when 4717 => read_data_o <= x"0000";
when 4718 => read_data_o <= x"0000";
when 4719 => read_data_o <= x"0000";
when 4720 => read_data_o <= x"0000";
when 4721 => read_data_o <= x"0000";
when 4722 => read_data_o <= x"0000";
when 4723 => read_data_o <= x"0000";
when 4724 => read_data_o <= x"0000";
when 4725 => read_data_o <= x"0000";
when 4726 => read_data_o <= x"0000";
when 4727 => read_data_o <= x"0000";
when 4728 => read_data_o <= x"0000";
when 4729 => read_data_o <= x"0000";
when 4730 => read_data_o <= x"0000";
when 4731 => read_data_o <= x"0000";
when 4732 => read_data_o <= x"0000";
when 4733 => read_data_o <= x"0000";
when 4734 => read_data_o <= x"0000";
when 4735 => read_data_o <= x"0000";
when 4736 => read_data_o <= x"0000";
when 4737 => read_data_o <= x"0000";
when 4738 => read_data_o <= x"0000";
when 4739 => read_data_o <= x"0000";
when 4740 => read_data_o <= x"0000";
when 4741 => read_data_o <= x"0000";
when 4742 => read_data_o <= x"0000";
when 4743 => read_data_o <= x"0000";
when 4744 => read_data_o <= x"0000";
when 4745 => read_data_o <= x"0000";
when 4746 => read_data_o <= x"0000";
when 4747 => read_data_o <= x"0000";
when 4748 => read_data_o <= x"0000";
when 4749 => read_data_o <= x"0000";
when 4750 => read_data_o <= x"0000";
when 4751 => read_data_o <= x"0000";
when 4752 => read_data_o <= x"0000";
when 4753 => read_data_o <= x"0000";
when 4754 => read_data_o <= x"0000";
when 4755 => read_data_o <= x"0000";
when 4756 => read_data_o <= x"0000";
when 4757 => read_data_o <= x"0000";
when 4758 => read_data_o <= x"0000";
when 4759 => read_data_o <= x"0000";
when 4760 => read_data_o <= x"0000";
when 4761 => read_data_o <= x"0000";
when 4762 => read_data_o <= x"0000";
when 4763 => read_data_o <= x"0000";
when 4764 => read_data_o <= x"0000";
when 4765 => read_data_o <= x"0000";
when 4766 => read_data_o <= x"0000";
when 4767 => read_data_o <= x"0000";
when 4768 => read_data_o <= x"0000";
when 4769 => read_data_o <= x"0000";
when 4770 => read_data_o <= x"0000";
when 4771 => read_data_o <= x"0000";
when 4772 => read_data_o <= x"d770";
when 4773 => read_data_o <= x"041a";
when 4774 => read_data_o <= x"0000";
when 4775 => read_data_o <= x"0000";
when 4776 => read_data_o <= x"0001";
when 4777 => read_data_o <= x"0000";
when 4778 => read_data_o <= x"0000";
when 4779 => read_data_o <= x"0000";
when 4780 => read_data_o <= x"0000";
when 4781 => read_data_o <= x"0000";
when 4782 => read_data_o <= x"0000";
when 4783 => read_data_o <= x"0000";
when 4784 => read_data_o <= x"0000";
when 4785 => read_data_o <= x"0000";
when 4786 => read_data_o <= x"0000";
when 4787 => read_data_o <= x"0000";
when 4788 => read_data_o <= x"0000";
when 4789 => read_data_o <= x"0000";
when 4790 => read_data_o <= x"0000";
when 4791 => read_data_o <= x"0000";
when 4792 => read_data_o <= x"0000";
when 4793 => read_data_o <= x"0000";
when 4794 => read_data_o <= x"0000";
when 4795 => read_data_o <= x"0000";
when 4796 => read_data_o <= x"0000";
when 4797 => read_data_o <= x"0000";
when 4798 => read_data_o <= x"0000";
when 4799 => read_data_o <= x"0000";
when 4800 => read_data_o <= x"0000";
when 4801 => read_data_o <= x"0000";
when 4802 => read_data_o <= x"0000";
when 4803 => read_data_o <= x"0000";
when 4804 => read_data_o <= x"0000";
when 4805 => read_data_o <= x"0000";
when 4806 => read_data_o <= x"0000";
when 4807 => read_data_o <= x"0000";
when 4808 => read_data_o <= x"0000";
when 4809 => read_data_o <= x"0000";
when 4810 => read_data_o <= x"0000";
when 4811 => read_data_o <= x"0000";
when 4812 => read_data_o <= x"0000";
when 4813 => read_data_o <= x"0000";
when 4814 => read_data_o <= x"0000";
when 4815 => read_data_o <= x"0000";
when 4816 => read_data_o <= x"0000";
when 4817 => read_data_o <= x"0000";
when 4818 => read_data_o <= x"0000";
when 4819 => read_data_o <= x"0000";
when 4820 => read_data_o <= x"0000";
when 4821 => read_data_o <= x"0000";
when 4822 => read_data_o <= x"0000";
when 4823 => read_data_o <= x"0000";
when 4824 => read_data_o <= x"0000";
when 4825 => read_data_o <= x"0000";
when 4826 => read_data_o <= x"0000";
when 4827 => read_data_o <= x"0000";
when 4828 => read_data_o <= x"0000";
when 4829 => read_data_o <= x"0000";
when 4830 => read_data_o <= x"0000";
when 4831 => read_data_o <= x"0000";
when 4832 => read_data_o <= x"0000";
when 4833 => read_data_o <= x"0000";
when 4834 => read_data_o <= x"0000";
when 4835 => read_data_o <= x"0000";
when 4836 => read_data_o <= x"0000";
when 4837 => read_data_o <= x"0000";
when 4838 => read_data_o <= x"0000";
when 4839 => read_data_o <= x"0000";
when 4840 => read_data_o <= x"0000";
when 4841 => read_data_o <= x"0000";
when 4842 => read_data_o <= x"0000";
when 4843 => read_data_o <= x"0000";
when 4844 => read_data_o <= x"0000";
when 4845 => read_data_o <= x"0000";
when 4846 => read_data_o <= x"0000";
when 4847 => read_data_o <= x"0000";
when 4848 => read_data_o <= x"0000";
when 4849 => read_data_o <= x"0000";
when 4850 => read_data_o <= x"0000";
when 4851 => read_data_o <= x"0000";
when 4852 => read_data_o <= x"d770";
when 4853 => read_data_o <= x"041a";
when 4854 => read_data_o <= x"0000";
when 4855 => read_data_o <= x"0000";
when 4856 => read_data_o <= x"0002";
when 4857 => read_data_o <= x"0000";
when 4858 => read_data_o <= x"0000";
when 4859 => read_data_o <= x"0000";
when 4860 => read_data_o <= x"0000";
when 4861 => read_data_o <= x"0000";
when 4862 => read_data_o <= x"0000";
when 4863 => read_data_o <= x"0000";
when 4864 => read_data_o <= x"0000";
when 4865 => read_data_o <= x"0000";
when 4866 => read_data_o <= x"0000";
when 4867 => read_data_o <= x"0000";
when 4868 => read_data_o <= x"0000";
when 4869 => read_data_o <= x"0000";
when 4870 => read_data_o <= x"0000";
when 4871 => read_data_o <= x"0000";
when 4872 => read_data_o <= x"0000";
when 4873 => read_data_o <= x"0000";
when 4874 => read_data_o <= x"0000";
when 4875 => read_data_o <= x"0000";
when 4876 => read_data_o <= x"0000";
when 4877 => read_data_o <= x"0000";
when 4878 => read_data_o <= x"0000";
when 4879 => read_data_o <= x"0000";
when 4880 => read_data_o <= x"0000";
when 4881 => read_data_o <= x"0000";
when 4882 => read_data_o <= x"0000";
when 4883 => read_data_o <= x"0000";
when 4884 => read_data_o <= x"0000";
when 4885 => read_data_o <= x"0000";
when 4886 => read_data_o <= x"0000";
when 4887 => read_data_o <= x"0000";
when 4888 => read_data_o <= x"0000";
when 4889 => read_data_o <= x"0000";
when 4890 => read_data_o <= x"0000";
when 4891 => read_data_o <= x"0000";
when 4892 => read_data_o <= x"0000";
when 4893 => read_data_o <= x"0000";
when 4894 => read_data_o <= x"0000";
when 4895 => read_data_o <= x"0000";
when 4896 => read_data_o <= x"0000";
when 4897 => read_data_o <= x"0000";
when 4898 => read_data_o <= x"0000";
when 4899 => read_data_o <= x"0000";
when 4900 => read_data_o <= x"0000";
when 4901 => read_data_o <= x"0000";
when 4902 => read_data_o <= x"0000";
when 4903 => read_data_o <= x"0000";
when 4904 => read_data_o <= x"0000";
when 4905 => read_data_o <= x"0000";
when 4906 => read_data_o <= x"0000";
when 4907 => read_data_o <= x"0000";
when 4908 => read_data_o <= x"0000";
when 4909 => read_data_o <= x"0000";
when 4910 => read_data_o <= x"0000";
when 4911 => read_data_o <= x"0000";
when 4912 => read_data_o <= x"0000";
when 4913 => read_data_o <= x"0000";
when 4914 => read_data_o <= x"0000";
when 4915 => read_data_o <= x"0000";
when 4916 => read_data_o <= x"0000";
when 4917 => read_data_o <= x"0000";
when 4918 => read_data_o <= x"0000";
when 4919 => read_data_o <= x"0000";
when 4920 => read_data_o <= x"0000";
when 4921 => read_data_o <= x"0000";
when 4922 => read_data_o <= x"0000";
when 4923 => read_data_o <= x"0000";
when 4924 => read_data_o <= x"0000";
when 4925 => read_data_o <= x"0000";
when 4926 => read_data_o <= x"0000";
when 4927 => read_data_o <= x"0000";
when 4928 => read_data_o <= x"0000";
when 4929 => read_data_o <= x"0000";
when 4930 => read_data_o <= x"7978";
when 4931 => read_data_o <= x"7400";
when 4932 => read_data_o <= x"d770";
when 4933 => read_data_o <= x"041a";
when 4934 => read_data_o <= x"0000";
when 4935 => read_data_o <= x"0000";
when 4936 => read_data_o <= x"0003";
when 4937 => read_data_o <= x"0000";
when 4938 => read_data_o <= x"0000";
when 4939 => read_data_o <= x"0000";
when 4940 => read_data_o <= x"0000";
when 4941 => read_data_o <= x"0000";
when 4942 => read_data_o <= x"0000";
when 4943 => read_data_o <= x"0000";
when 4944 => read_data_o <= x"0000";
when 4945 => read_data_o <= x"0000";
when 4946 => read_data_o <= x"0000";
when 4947 => read_data_o <= x"0000";
when 4948 => read_data_o <= x"0000";
when 4949 => read_data_o <= x"0000";
when 4950 => read_data_o <= x"0000";
when 4951 => read_data_o <= x"0000";
when 4952 => read_data_o <= x"0000";
when 4953 => read_data_o <= x"0000";
when 4954 => read_data_o <= x"0000";
when 4955 => read_data_o <= x"0000";
when 4956 => read_data_o <= x"0000";
when 4957 => read_data_o <= x"0000";
when 4958 => read_data_o <= x"0000";
when 4959 => read_data_o <= x"0000";
when 4960 => read_data_o <= x"0000";
when 4961 => read_data_o <= x"0000";
when 4962 => read_data_o <= x"0000";
when 4963 => read_data_o <= x"0000";
when 4964 => read_data_o <= x"0000";
when 4965 => read_data_o <= x"0000";
when 4966 => read_data_o <= x"0000";
when 4967 => read_data_o <= x"0000";
when 4968 => read_data_o <= x"0000";
when 4969 => read_data_o <= x"0000";
when 4970 => read_data_o <= x"0000";
when 4971 => read_data_o <= x"0000";
when 4972 => read_data_o <= x"0000";
when 4973 => read_data_o <= x"0000";
when 4974 => read_data_o <= x"0000";
when 4975 => read_data_o <= x"0000";
when 4976 => read_data_o <= x"0000";
when 4977 => read_data_o <= x"0000";
when 4978 => read_data_o <= x"0000";
when 4979 => read_data_o <= x"0000";
when 4980 => read_data_o <= x"0000";
when 4981 => read_data_o <= x"0000";
when 4982 => read_data_o <= x"0000";
when 4983 => read_data_o <= x"0000";
when 4984 => read_data_o <= x"0000";
when 4985 => read_data_o <= x"0000";
when 4986 => read_data_o <= x"0000";
when 4987 => read_data_o <= x"0000";
when 4988 => read_data_o <= x"0000";
when 4989 => read_data_o <= x"0000";
when 4990 => read_data_o <= x"0000";
when 4991 => read_data_o <= x"0000";
when 4992 => read_data_o <= x"0000";
when 4993 => read_data_o <= x"0000";
when 4994 => read_data_o <= x"0000";
when 4995 => read_data_o <= x"0000";
when 4996 => read_data_o <= x"0000";
when 4997 => read_data_o <= x"0000";
when 4998 => read_data_o <= x"0000";
when 4999 => read_data_o <= x"0000";
when 5000 => read_data_o <= x"0000";
when 5001 => read_data_o <= x"0000";
when 5002 => read_data_o <= x"0000";
when 5003 => read_data_o <= x"0000";
when 5004 => read_data_o <= x"0000";
when 5005 => read_data_o <= x"0000";
when 5006 => read_data_o <= x"0000";
when 5007 => read_data_o <= x"0000";
when 5008 => read_data_o <= x"0000";
when 5009 => read_data_o <= x"0000";
when 5010 => read_data_o <= x"0000";
when 5011 => read_data_o <= x"0000";
when 5012 => read_data_o <= x"d770";
when 5013 => read_data_o <= x"041a";
when 5014 => read_data_o <= x"0000";
when 5015 => read_data_o <= x"0000";
when 5016 => read_data_o <= x"0004";
when 5017 => read_data_o <= x"0000";
when 5018 => read_data_o <= x"0000";
when 5019 => read_data_o <= x"0000";
when 5020 => read_data_o <= x"0000";
when 5021 => read_data_o <= x"0000";
when 5022 => read_data_o <= x"0000";
when 5023 => read_data_o <= x"0000";
when 5024 => read_data_o <= x"0000";
when 5025 => read_data_o <= x"0000";
when 5026 => read_data_o <= x"0000";
when 5027 => read_data_o <= x"0000";
when 5028 => read_data_o <= x"0000";
when 5029 => read_data_o <= x"0000";
when 5030 => read_data_o <= x"0000";
when 5031 => read_data_o <= x"0000";
when 5032 => read_data_o <= x"0000";
when 5033 => read_data_o <= x"0000";
when 5034 => read_data_o <= x"0000";
when 5035 => read_data_o <= x"0000";
when 5036 => read_data_o <= x"0000";
when 5037 => read_data_o <= x"0000";
when 5038 => read_data_o <= x"0000";
when 5039 => read_data_o <= x"0000";
when 5040 => read_data_o <= x"0000";
when 5041 => read_data_o <= x"0000";
when 5042 => read_data_o <= x"0000";
when 5043 => read_data_o <= x"0000";
when 5044 => read_data_o <= x"0000";
when 5045 => read_data_o <= x"0000";
when 5046 => read_data_o <= x"0000";
when 5047 => read_data_o <= x"0000";
when 5048 => read_data_o <= x"0000";
when 5049 => read_data_o <= x"0000";
when 5050 => read_data_o <= x"0000";
when 5051 => read_data_o <= x"0000";
when 5052 => read_data_o <= x"0000";
when 5053 => read_data_o <= x"0000";
when 5054 => read_data_o <= x"0000";
when 5055 => read_data_o <= x"0000";
when 5056 => read_data_o <= x"0000";
when 5057 => read_data_o <= x"0000";
when 5058 => read_data_o <= x"0000";
when 5059 => read_data_o <= x"0000";
when 5060 => read_data_o <= x"0000";
when 5061 => read_data_o <= x"0000";
when 5062 => read_data_o <= x"0000";
when 5063 => read_data_o <= x"0000";
when 5064 => read_data_o <= x"0000";
when 5065 => read_data_o <= x"0000";
when 5066 => read_data_o <= x"0000";
when 5067 => read_data_o <= x"0000";
when 5068 => read_data_o <= x"0000";
when 5069 => read_data_o <= x"0000";
when 5070 => read_data_o <= x"0000";
when 5071 => read_data_o <= x"0000";
when 5072 => read_data_o <= x"0000";
when 5073 => read_data_o <= x"0000";
when 5074 => read_data_o <= x"0000";
when 5075 => read_data_o <= x"0000";
when 5076 => read_data_o <= x"0000";
when 5077 => read_data_o <= x"0000";
when 5078 => read_data_o <= x"0000";
when 5079 => read_data_o <= x"0000";
when 5080 => read_data_o <= x"0000";
when 5081 => read_data_o <= x"0000";
when 5082 => read_data_o <= x"0000";
when 5083 => read_data_o <= x"0000";
when 5084 => read_data_o <= x"0000";
when 5085 => read_data_o <= x"0000";
when 5086 => read_data_o <= x"0000";
when 5087 => read_data_o <= x"0000";
when 5088 => read_data_o <= x"0000";
when 5089 => read_data_o <= x"0000";
when 5090 => read_data_o <= x"0000";
when 5091 => read_data_o <= x"0000";
when 5092 => read_data_o <= x"d770";
when 5093 => read_data_o <= x"041a";
when 5094 => read_data_o <= x"0000";
when 5095 => read_data_o <= x"0000";
when 5096 => read_data_o <= x"0005";
when 5097 => read_data_o <= x"0000";
when 5098 => read_data_o <= x"0000";
when 5099 => read_data_o <= x"0000";
when 5100 => read_data_o <= x"0000";
when 5101 => read_data_o <= x"0000";
when 5102 => read_data_o <= x"0000";
when 5103 => read_data_o <= x"0000";
when 5104 => read_data_o <= x"0000";
when 5105 => read_data_o <= x"0000";
when 5106 => read_data_o <= x"0000";
when 5107 => read_data_o <= x"0000";
when 5108 => read_data_o <= x"0000";
when 5109 => read_data_o <= x"0000";
when 5110 => read_data_o <= x"0000";
when 5111 => read_data_o <= x"0000";
when 5112 => read_data_o <= x"0000";
when 5113 => read_data_o <= x"0000";
when 5114 => read_data_o <= x"0000";
when 5115 => read_data_o <= x"0000";
when 5116 => read_data_o <= x"0000";
when 5117 => read_data_o <= x"0000";
when 5118 => read_data_o <= x"0000";
when 5119 => read_data_o <= x"0000";
when 5120 => read_data_o <= x"0000";
when 5121 => read_data_o <= x"0000";
when 5122 => read_data_o <= x"0000";
when 5123 => read_data_o <= x"0000";
when 5124 => read_data_o <= x"0000";
when 5125 => read_data_o <= x"0000";
when 5126 => read_data_o <= x"0000";
when 5127 => read_data_o <= x"0000";
when 5128 => read_data_o <= x"0000";
when 5129 => read_data_o <= x"0000";
when 5130 => read_data_o <= x"0000";
when 5131 => read_data_o <= x"0000";
when 5132 => read_data_o <= x"0000";
when 5133 => read_data_o <= x"0000";
when 5134 => read_data_o <= x"0000";
when 5135 => read_data_o <= x"0000";
when 5136 => read_data_o <= x"0000";
when 5137 => read_data_o <= x"0000";
when 5138 => read_data_o <= x"0000";
when 5139 => read_data_o <= x"0000";
when 5140 => read_data_o <= x"0000";
when 5141 => read_data_o <= x"0000";
when 5142 => read_data_o <= x"0000";
when 5143 => read_data_o <= x"0000";
when 5144 => read_data_o <= x"0000";
when 5145 => read_data_o <= x"0000";
when 5146 => read_data_o <= x"0000";
when 5147 => read_data_o <= x"0000";
when 5148 => read_data_o <= x"0000";
when 5149 => read_data_o <= x"0000";
when 5150 => read_data_o <= x"0000";
when 5151 => read_data_o <= x"0000";
when 5152 => read_data_o <= x"0000";
when 5153 => read_data_o <= x"0000";
when 5154 => read_data_o <= x"0000";
when 5155 => read_data_o <= x"0000";
when 5156 => read_data_o <= x"0000";
when 5157 => read_data_o <= x"0000";
when 5158 => read_data_o <= x"0000";
when 5159 => read_data_o <= x"0000";
when 5160 => read_data_o <= x"0000";
when 5161 => read_data_o <= x"0000";
when 5162 => read_data_o <= x"0000";
when 5163 => read_data_o <= x"0000";
when 5164 => read_data_o <= x"0000";
when 5165 => read_data_o <= x"0000";
when 5166 => read_data_o <= x"0000";
when 5167 => read_data_o <= x"0000";
when 5168 => read_data_o <= x"0000";
when 5169 => read_data_o <= x"0000";
when 5170 => read_data_o <= x"0000";
when 5171 => read_data_o <= x"0000";
when 5172 => read_data_o <= x"d770";
when 5173 => read_data_o <= x"041a";
when 5174 => read_data_o <= x"0000";
when 5175 => read_data_o <= x"0000";
when 5176 => read_data_o <= x"0006";
when 5177 => read_data_o <= x"0000";
when 5178 => read_data_o <= x"0000";
when 5179 => read_data_o <= x"0000";
when 5180 => read_data_o <= x"0000";
when 5181 => read_data_o <= x"0000";
when 5182 => read_data_o <= x"0000";
when 5183 => read_data_o <= x"0000";
when 5184 => read_data_o <= x"0000";
when 5185 => read_data_o <= x"0000";
when 5186 => read_data_o <= x"0000";
when 5187 => read_data_o <= x"0000";
when 5188 => read_data_o <= x"0000";
when 5189 => read_data_o <= x"0000";
when 5190 => read_data_o <= x"0000";
when 5191 => read_data_o <= x"0000";
when 5192 => read_data_o <= x"0000";
when 5193 => read_data_o <= x"0000";
when 5194 => read_data_o <= x"0000";
when 5195 => read_data_o <= x"0000";
when 5196 => read_data_o <= x"0000";
when 5197 => read_data_o <= x"0000";
when 5198 => read_data_o <= x"0000";
when 5199 => read_data_o <= x"0000";
when 5200 => read_data_o <= x"0000";
when 5201 => read_data_o <= x"0000";
when 5202 => read_data_o <= x"0000";
when 5203 => read_data_o <= x"0000";
when 5204 => read_data_o <= x"0000";
when 5205 => read_data_o <= x"0000";
when 5206 => read_data_o <= x"0000";
when 5207 => read_data_o <= x"0000";
when 5208 => read_data_o <= x"0000";
when 5209 => read_data_o <= x"0000";
when 5210 => read_data_o <= x"0000";
when 5211 => read_data_o <= x"0000";
when 5212 => read_data_o <= x"0000";
when 5213 => read_data_o <= x"0000";
when 5214 => read_data_o <= x"0000";
when 5215 => read_data_o <= x"0000";
when 5216 => read_data_o <= x"0000";
when 5217 => read_data_o <= x"0000";
when 5218 => read_data_o <= x"0000";
when 5219 => read_data_o <= x"0000";
when 5220 => read_data_o <= x"0000";
when 5221 => read_data_o <= x"0000";
when 5222 => read_data_o <= x"0000";
when 5223 => read_data_o <= x"0000";
when 5224 => read_data_o <= x"0000";
when 5225 => read_data_o <= x"0000";
when 5226 => read_data_o <= x"0000";
when 5227 => read_data_o <= x"0000";
when 5228 => read_data_o <= x"0000";
when 5229 => read_data_o <= x"0000";
when 5230 => read_data_o <= x"0000";
when 5231 => read_data_o <= x"0000";
when 5232 => read_data_o <= x"0000";
when 5233 => read_data_o <= x"0000";
when 5234 => read_data_o <= x"0000";
when 5235 => read_data_o <= x"0000";
when 5236 => read_data_o <= x"0000";
when 5237 => read_data_o <= x"0000";
when 5238 => read_data_o <= x"0000";
when 5239 => read_data_o <= x"0000";
when 5240 => read_data_o <= x"0000";
when 5241 => read_data_o <= x"0000";
when 5242 => read_data_o <= x"0000";
when 5243 => read_data_o <= x"0000";
when 5244 => read_data_o <= x"0000";
when 5245 => read_data_o <= x"0000";
when 5246 => read_data_o <= x"0000";
when 5247 => read_data_o <= x"0000";
when 5248 => read_data_o <= x"0000";
when 5249 => read_data_o <= x"0000";
when 5250 => read_data_o <= x"0073";
when 5251 => read_data_o <= x"6576";
when 5252 => read_data_o <= x"d770";
when 5253 => read_data_o <= x"041a";
when 5254 => read_data_o <= x"0000";
when 5255 => read_data_o <= x"0000";
when 5256 => read_data_o <= x"0007";
when 5257 => read_data_o <= x"0000";
when 5258 => read_data_o <= x"0000";
when 5259 => read_data_o <= x"0000";
when 5260 => read_data_o <= x"0000";
when 5261 => read_data_o <= x"0000";
when 5262 => read_data_o <= x"0000";
when 5263 => read_data_o <= x"0000";
when 5264 => read_data_o <= x"0000";
when 5265 => read_data_o <= x"0000";
when 5266 => read_data_o <= x"0000";
when 5267 => read_data_o <= x"0000";
when 5268 => read_data_o <= x"0000";
when 5269 => read_data_o <= x"0000";
when 5270 => read_data_o <= x"0000";
when 5271 => read_data_o <= x"0000";
when 5272 => read_data_o <= x"0000";
when 5273 => read_data_o <= x"0000";
when 5274 => read_data_o <= x"0000";
when 5275 => read_data_o <= x"0000";
when 5276 => read_data_o <= x"0000";
when 5277 => read_data_o <= x"0000";
when 5278 => read_data_o <= x"0000";
when 5279 => read_data_o <= x"0000";
when 5280 => read_data_o <= x"0000";
when 5281 => read_data_o <= x"0000";
when 5282 => read_data_o <= x"0000";
when 5283 => read_data_o <= x"0000";
when 5284 => read_data_o <= x"0000";
when 5285 => read_data_o <= x"0000";
when 5286 => read_data_o <= x"0000";
when 5287 => read_data_o <= x"0000";
when 5288 => read_data_o <= x"0000";
when 5289 => read_data_o <= x"0000";
when 5290 => read_data_o <= x"0000";
when 5291 => read_data_o <= x"0000";
when 5292 => read_data_o <= x"0000";
when 5293 => read_data_o <= x"0000";
when 5294 => read_data_o <= x"0000";
when 5295 => read_data_o <= x"0000";
when 5296 => read_data_o <= x"0000";
when 5297 => read_data_o <= x"0000";
when 5298 => read_data_o <= x"0000";
when 5299 => read_data_o <= x"0000";
when 5300 => read_data_o <= x"0000";
when 5301 => read_data_o <= x"0000";
when 5302 => read_data_o <= x"0000";
when 5303 => read_data_o <= x"0000";
when 5304 => read_data_o <= x"0000";
when 5305 => read_data_o <= x"0000";
when 5306 => read_data_o <= x"0000";
when 5307 => read_data_o <= x"0000";
when 5308 => read_data_o <= x"0000";
when 5309 => read_data_o <= x"0000";
when 5310 => read_data_o <= x"0000";
when 5311 => read_data_o <= x"0000";
when 5312 => read_data_o <= x"0000";
when 5313 => read_data_o <= x"0000";
when 5314 => read_data_o <= x"0000";
when 5315 => read_data_o <= x"0000";
when 5316 => read_data_o <= x"0000";
when 5317 => read_data_o <= x"0000";
when 5318 => read_data_o <= x"0000";
when 5319 => read_data_o <= x"0000";
when 5320 => read_data_o <= x"0000";
when 5321 => read_data_o <= x"0000";
when 5322 => read_data_o <= x"0000";
when 5323 => read_data_o <= x"0000";
when 5324 => read_data_o <= x"0000";
when 5325 => read_data_o <= x"0000";
when 5326 => read_data_o <= x"0000";
when 5327 => read_data_o <= x"0000";
when 5328 => read_data_o <= x"0000";
when 5329 => read_data_o <= x"0000";
when 5330 => read_data_o <= x"0000";
when 5331 => read_data_o <= x"0000";
when 5332 => read_data_o <= x"d770";
when 5333 => read_data_o <= x"041a";
when 5334 => read_data_o <= x"0000";
when 5335 => read_data_o <= x"0000";
when 5336 => read_data_o <= x"0008";
when 5337 => read_data_o <= x"0000";
when 5338 => read_data_o <= x"0000";
when 5339 => read_data_o <= x"0000";
when 5340 => read_data_o <= x"0000";
when 5341 => read_data_o <= x"0000";
when 5342 => read_data_o <= x"0000";
when 5343 => read_data_o <= x"0000";
when 5344 => read_data_o <= x"0000";
when 5345 => read_data_o <= x"0000";
when 5346 => read_data_o <= x"0000";
when 5347 => read_data_o <= x"0000";
when 5348 => read_data_o <= x"0000";
when 5349 => read_data_o <= x"0000";
when 5350 => read_data_o <= x"0000";
when 5351 => read_data_o <= x"0000";
when 5352 => read_data_o <= x"0000";
when 5353 => read_data_o <= x"0000";
when 5354 => read_data_o <= x"0000";
when 5355 => read_data_o <= x"0000";
when 5356 => read_data_o <= x"0000";
when 5357 => read_data_o <= x"0000";
when 5358 => read_data_o <= x"0000";
when 5359 => read_data_o <= x"0000";
when 5360 => read_data_o <= x"0000";
when 5361 => read_data_o <= x"0000";
when 5362 => read_data_o <= x"0000";
when 5363 => read_data_o <= x"0000";
when 5364 => read_data_o <= x"0000";
when 5365 => read_data_o <= x"0000";
when 5366 => read_data_o <= x"0000";
when 5367 => read_data_o <= x"0000";
when 5368 => read_data_o <= x"0000";
when 5369 => read_data_o <= x"0000";
when 5370 => read_data_o <= x"0000";
when 5371 => read_data_o <= x"0000";
when 5372 => read_data_o <= x"0000";
when 5373 => read_data_o <= x"0000";
when 5374 => read_data_o <= x"0000";
when 5375 => read_data_o <= x"0000";
when 5376 => read_data_o <= x"0000";
when 5377 => read_data_o <= x"0000";
when 5378 => read_data_o <= x"0000";
when 5379 => read_data_o <= x"0000";
when 5380 => read_data_o <= x"0000";
when 5381 => read_data_o <= x"0000";
when 5382 => read_data_o <= x"0000";
when 5383 => read_data_o <= x"0000";
when 5384 => read_data_o <= x"0000";
when 5385 => read_data_o <= x"0000";
when 5386 => read_data_o <= x"0000";
when 5387 => read_data_o <= x"0000";
when 5388 => read_data_o <= x"0000";
when 5389 => read_data_o <= x"0000";
when 5390 => read_data_o <= x"0000";
when 5391 => read_data_o <= x"0000";
when 5392 => read_data_o <= x"0000";
when 5393 => read_data_o <= x"0000";
when 5394 => read_data_o <= x"0000";
when 5395 => read_data_o <= x"0000";
when 5396 => read_data_o <= x"0000";
when 5397 => read_data_o <= x"0000";
when 5398 => read_data_o <= x"0000";
when 5399 => read_data_o <= x"0000";
when 5400 => read_data_o <= x"0000";
when 5401 => read_data_o <= x"0000";
when 5402 => read_data_o <= x"0000";
when 5403 => read_data_o <= x"0000";
when 5404 => read_data_o <= x"0000";
when 5405 => read_data_o <= x"0000";
when 5406 => read_data_o <= x"0000";
when 5407 => read_data_o <= x"0000";
when 5408 => read_data_o <= x"0000";
when 5409 => read_data_o <= x"0000";
when 5410 => read_data_o <= x"0000";
when 5411 => read_data_o <= x"0000";
when 5412 => read_data_o <= x"d770";
when 5413 => read_data_o <= x"041a";
when 5414 => read_data_o <= x"0000";
when 5415 => read_data_o <= x"0000";
when 5416 => read_data_o <= x"0009";
when 5417 => read_data_o <= x"0000";
when 5418 => read_data_o <= x"0000";
when 5419 => read_data_o <= x"0000";
when 5420 => read_data_o <= x"0000";
when 5421 => read_data_o <= x"0000";
when 5422 => read_data_o <= x"0000";
when 5423 => read_data_o <= x"0000";
when 5424 => read_data_o <= x"0000";
when 5425 => read_data_o <= x"0000";
when 5426 => read_data_o <= x"0000";
when 5427 => read_data_o <= x"0000";
when 5428 => read_data_o <= x"0000";
when 5429 => read_data_o <= x"0000";
when 5430 => read_data_o <= x"0000";
when 5431 => read_data_o <= x"0000";
when 5432 => read_data_o <= x"0000";
when 5433 => read_data_o <= x"0000";
when 5434 => read_data_o <= x"0000";
when 5435 => read_data_o <= x"0000";
when 5436 => read_data_o <= x"0000";
when 5437 => read_data_o <= x"0000";
when 5438 => read_data_o <= x"0000";
when 5439 => read_data_o <= x"0000";
when 5440 => read_data_o <= x"0000";
when 5441 => read_data_o <= x"0000";
when 5442 => read_data_o <= x"0000";
when 5443 => read_data_o <= x"0000";
when 5444 => read_data_o <= x"0000";
when 5445 => read_data_o <= x"0000";
when 5446 => read_data_o <= x"0000";
when 5447 => read_data_o <= x"0000";
when 5448 => read_data_o <= x"0000";
when 5449 => read_data_o <= x"0000";
when 5450 => read_data_o <= x"0000";
when 5451 => read_data_o <= x"0000";
when 5452 => read_data_o <= x"0000";
when 5453 => read_data_o <= x"0000";
when 5454 => read_data_o <= x"0000";
when 5455 => read_data_o <= x"0000";
when 5456 => read_data_o <= x"0000";
when 5457 => read_data_o <= x"0000";
when 5458 => read_data_o <= x"0000";
when 5459 => read_data_o <= x"0000";
when 5460 => read_data_o <= x"0000";
when 5461 => read_data_o <= x"0000";
when 5462 => read_data_o <= x"0000";
when 5463 => read_data_o <= x"0000";
when 5464 => read_data_o <= x"0000";
when 5465 => read_data_o <= x"0000";
when 5466 => read_data_o <= x"0000";
when 5467 => read_data_o <= x"0000";
when 5468 => read_data_o <= x"0000";
when 5469 => read_data_o <= x"0000";
when 5470 => read_data_o <= x"0000";
when 5471 => read_data_o <= x"0000";
when 5472 => read_data_o <= x"0000";
when 5473 => read_data_o <= x"0000";
when 5474 => read_data_o <= x"0000";
when 5475 => read_data_o <= x"0000";
when 5476 => read_data_o <= x"0000";
when 5477 => read_data_o <= x"0000";
when 5478 => read_data_o <= x"0000";
when 5479 => read_data_o <= x"0000";
when 5480 => read_data_o <= x"0000";
when 5481 => read_data_o <= x"0000";
when 5482 => read_data_o <= x"0000";
when 5483 => read_data_o <= x"0000";
when 5484 => read_data_o <= x"0000";
when 5485 => read_data_o <= x"0000";
when 5486 => read_data_o <= x"0000";
when 5487 => read_data_o <= x"0000";
when 5488 => read_data_o <= x"0000";
when 5489 => read_data_o <= x"0000";
when 5490 => read_data_o <= x"0000";
when 5491 => read_data_o <= x"0000";
when 5492 => read_data_o <= x"d770";
when 5493 => read_data_o <= x"041a";
when 5494 => read_data_o <= x"0000";
when 5495 => read_data_o <= x"0000";
when 5496 => read_data_o <= x"000a";
when 5497 => read_data_o <= x"0000";
when 5498 => read_data_o <= x"0000";
when 5499 => read_data_o <= x"0000";
when 5500 => read_data_o <= x"0000";
when 5501 => read_data_o <= x"0000";
when 5502 => read_data_o <= x"0000";
when 5503 => read_data_o <= x"0079";
when 5504 => read_data_o <= x"0000";
when 5505 => read_data_o <= x"0000";
when 5506 => read_data_o <= x"0000";
when 5507 => read_data_o <= x"0000";
when 5508 => read_data_o <= x"0000";
when 5509 => read_data_o <= x"0000";
when 5510 => read_data_o <= x"0000";
when 5511 => read_data_o <= x"0000";
when 5512 => read_data_o <= x"0000";
when 5513 => read_data_o <= x"0000";
when 5514 => read_data_o <= x"0000";
when 5515 => read_data_o <= x"0000";
when 5516 => read_data_o <= x"0000";
when 5517 => read_data_o <= x"0000";
when 5518 => read_data_o <= x"0000";
when 5519 => read_data_o <= x"0000";
when 5520 => read_data_o <= x"0000";
when 5521 => read_data_o <= x"0000";
when 5522 => read_data_o <= x"0000";
when 5523 => read_data_o <= x"0000";
when 5524 => read_data_o <= x"0000";
when 5525 => read_data_o <= x"0000";
when 5526 => read_data_o <= x"0000";
when 5527 => read_data_o <= x"0000";
when 5528 => read_data_o <= x"0000";
when 5529 => read_data_o <= x"0000";
when 5530 => read_data_o <= x"0000";
when 5531 => read_data_o <= x"0000";
when 5532 => read_data_o <= x"0000";
when 5533 => read_data_o <= x"0000";
when 5534 => read_data_o <= x"0000";
when 5535 => read_data_o <= x"0000";
when 5536 => read_data_o <= x"0000";
when 5537 => read_data_o <= x"0000";
when 5538 => read_data_o <= x"0000";
when 5539 => read_data_o <= x"0000";
when 5540 => read_data_o <= x"0000";
when 5541 => read_data_o <= x"0000";
when 5542 => read_data_o <= x"0000";
when 5543 => read_data_o <= x"0000";
when 5544 => read_data_o <= x"0000";
when 5545 => read_data_o <= x"0000";
when 5546 => read_data_o <= x"0000";
when 5547 => read_data_o <= x"0000";
when 5548 => read_data_o <= x"0000";
when 5549 => read_data_o <= x"0000";
when 5550 => read_data_o <= x"0000";
when 5551 => read_data_o <= x"0000";
when 5552 => read_data_o <= x"0000";
when 5553 => read_data_o <= x"0000";
when 5554 => read_data_o <= x"0000";
when 5555 => read_data_o <= x"0000";
when 5556 => read_data_o <= x"0000";
when 5557 => read_data_o <= x"0000";
when 5558 => read_data_o <= x"0000";
when 5559 => read_data_o <= x"0000";
when 5560 => read_data_o <= x"0000";
when 5561 => read_data_o <= x"0000";
when 5562 => read_data_o <= x"0000";
when 5563 => read_data_o <= x"0000";
when 5564 => read_data_o <= x"0000";
when 5565 => read_data_o <= x"0000";
when 5566 => read_data_o <= x"0000";
when 5567 => read_data_o <= x"0000";
when 5568 => read_data_o <= x"0000";
when 5569 => read_data_o <= x"0000";
when 5570 => read_data_o <= x"0000";
when 5571 => read_data_o <= x"0000";
when 5572 => read_data_o <= x"d770";
when 5573 => read_data_o <= x"041a";
when 5574 => read_data_o <= x"0000";
when 5575 => read_data_o <= x"0000";
when 5576 => read_data_o <= x"000b";
when 5577 => read_data_o <= x"0000";
when 5578 => read_data_o <= x"0000";
when 5579 => read_data_o <= x"0000";
when 5580 => read_data_o <= x"0000";
when 5581 => read_data_o <= x"0000";
when 5582 => read_data_o <= x"0000";
when 5583 => read_data_o <= x"0000";
when 5584 => read_data_o <= x"0000";
when 5585 => read_data_o <= x"0000";
when 5586 => read_data_o <= x"0000";
when 5587 => read_data_o <= x"0000";
when 5588 => read_data_o <= x"0000";
when 5589 => read_data_o <= x"0000";
when 5590 => read_data_o <= x"0000";
when 5591 => read_data_o <= x"0000";
when 5592 => read_data_o <= x"0000";
when 5593 => read_data_o <= x"0000";
when 5594 => read_data_o <= x"0000";
when 5595 => read_data_o <= x"0000";
when 5596 => read_data_o <= x"0000";
when 5597 => read_data_o <= x"0000";
when 5598 => read_data_o <= x"0000";
when 5599 => read_data_o <= x"0000";
when 5600 => read_data_o <= x"0000";
when 5601 => read_data_o <= x"0000";
when 5602 => read_data_o <= x"0000";
when 5603 => read_data_o <= x"0000";
when 5604 => read_data_o <= x"0000";
when 5605 => read_data_o <= x"0000";
when 5606 => read_data_o <= x"0000";
when 5607 => read_data_o <= x"0000";
when 5608 => read_data_o <= x"0000";
when 5609 => read_data_o <= x"0000";
when 5610 => read_data_o <= x"0000";
when 5611 => read_data_o <= x"0000";
when 5612 => read_data_o <= x"0000";
when 5613 => read_data_o <= x"0000";
when 5614 => read_data_o <= x"0000";
when 5615 => read_data_o <= x"0000";
when 5616 => read_data_o <= x"0000";
when 5617 => read_data_o <= x"0000";
when 5618 => read_data_o <= x"0000";
when 5619 => read_data_o <= x"0000";
when 5620 => read_data_o <= x"0000";
when 5621 => read_data_o <= x"0000";
when 5622 => read_data_o <= x"0000";
when 5623 => read_data_o <= x"0000";
when 5624 => read_data_o <= x"0000";
when 5625 => read_data_o <= x"0303";
when 5626 => read_data_o <= x"c2c2";
when 5627 => read_data_o <= x"8080";
when 5628 => read_data_o <= x"0000";
when 5629 => read_data_o <= x"0000";
when 5630 => read_data_o <= x"0000";
when 5631 => read_data_o <= x"0606";
when 5632 => read_data_o <= x"8585";
when 5633 => read_data_o <= x"0000";
when 5634 => read_data_o <= x"0000";
when 5635 => read_data_o <= x"0000";
when 5636 => read_data_o <= x"0000";
when 5637 => read_data_o <= x"0606";
when 5638 => read_data_o <= x"8585";
when 5639 => read_data_o <= x"0000";
when 5640 => read_data_o <= x"0000";
when 5641 => read_data_o <= x"f3f3";
when 5642 => read_data_o <= x"8080";
when 5643 => read_data_o <= x"0000";
when 5644 => read_data_o <= x"0000";
when 5645 => read_data_o <= x"0000";
when 5646 => read_data_o <= x"0000";
when 5647 => read_data_o <= x"0000";
when 5648 => read_data_o <= x"0000";
when 5649 => read_data_o <= x"0000";
when 5650 => read_data_o <= x"0808";
when 5651 => read_data_o <= x"5050";
when 5652 => read_data_o <= x"e8e8";
when 5653 => read_data_o <= x"0f0f";
when 5654 => read_data_o <= x"4040";
when 5655 => read_data_o <= x"0f0f";
when 5656 => read_data_o <= x"4040";
when 5657 => read_data_o <= x"0000";
when 5658 => read_data_o <= x"0000";
when 5659 => read_data_o <= x"e8e8";
when 5660 => read_data_o <= x"1818";
when 5661 => read_data_o <= x"0000";
when 5662 => read_data_o <= x"0000";
when 5663 => read_data_o <= x"0000";
when 5664 => read_data_o <= x"5050";
when 5665 => read_data_o <= x"0000";
when 5666 => read_data_o <= x"1010";
when 5667 => read_data_o <= x"5252";
when 5668 => read_data_o <= x"0000";
when 5669 => read_data_o <= x"6464";
when 5670 => read_data_o <= x"0000";
when 5671 => read_data_o <= x"0101";
when 5672 => read_data_o <= x"0000";
when 5673 => read_data_o <= x"0000";
when 5674 => read_data_o <= x"0101";
when 5675 => read_data_o <= x"0101";
when 5676 => read_data_o <= x"0000";
when 5677 => read_data_o <= x"0000";
when 5678 => read_data_o <= x"0202";
when 5679 => read_data_o <= x"8080";
when 5680 => read_data_o <= x"0000";
when 5681 => read_data_o <= x"0000";
when 5682 => read_data_o <= x"0303";
when 5683 => read_data_o <= x"0000";
when 5684 => read_data_o <= x"ffff";
when 5685 => read_data_o <= x"0101";
when 5686 => read_data_o <= x"2c2c";
when 5687 => read_data_o <= x"2c2c";
when 5688 => read_data_o <= x"2c2c";
when 5689 => read_data_o <= x"2c2c";
when 5690 => read_data_o <= x"2c2c";
when 5691 => read_data_o <= x"6464";
when 5692 => read_data_o <= x"6464";
when 5693 => read_data_o <= x"6464";
when 5694 => read_data_o <= x"6464";
when 5695 => read_data_o <= x"6464";
when 5696 => read_data_o <= x"5858";
when 5697 => read_data_o <= x"3838";
when 5698 => read_data_o <= x"d8d8";
when 5699 => read_data_o <= x"6464";
when 5700 => read_data_o <= x"0b0b";
when 5701 => read_data_o <= x"e8e8";
when 5702 => read_data_o <= x"0000";
when 5703 => read_data_o <= x"0000";
when 5704 => read_data_o <= x"0000";
when 5705 => read_data_o <= x"0000";
when 5706 => read_data_o <= x"0000";
when 5707 => read_data_o <= x"0000";
when 5708 => read_data_o <= x"0000";
when 5709 => read_data_o <= x"0000";
when 5710 => read_data_o <= x"ffff";
when 5711 => read_data_o <= x"2020";
when 5712 => read_data_o <= x"2020";
when 5713 => read_data_o <= x"2020";
when 5714 => read_data_o <= x"2020";
when 5715 => read_data_o <= x"2020";
when 5716 => read_data_o <= x"2020";
when 5717 => read_data_o <= x"5252";
when 5718 => read_data_o <= x"4545";
when 5719 => read_data_o <= x"0000";
when 5720 => read_data_o <= x"f0f0";
when 5721 => read_data_o <= x"f0f0";
when 5722 => read_data_o <= x"f0f0";
when 5723 => read_data_o <= x"f0f0";
when 5724 => read_data_o <= x"f0f0";
when 5725 => read_data_o <= x"0202";
when 5726 => read_data_o <= x"9b9b";
when 5727 => read_data_o <= x"c0c0";
when 5728 => read_data_o <= x"0202";
when 5729 => read_data_o <= x"9b9b";
when 5730 => read_data_o <= x"c0c0";
when 5731 => read_data_o <= x"0202";
when 5732 => read_data_o <= x"9b9b";
when 5733 => read_data_o <= x"c0c0";
when 5734 => read_data_o <= x"0202";
when 5735 => read_data_o <= x"9b9b";
when 5736 => read_data_o <= x"c0c0";
when 5737 => read_data_o <= x"0202";
when 5738 => read_data_o <= x"9b9b";
when 5739 => read_data_o <= x"c0c0";
when 5740 => read_data_o <= x"ffff";
when 5741 => read_data_o <= x"ffff";
when 5742 => read_data_o <= x"0a0a";
when 5743 => read_data_o <= x"0000";
when 5744 => read_data_o <= x"2020";
when 5745 => read_data_o <= x"2020";
when 5746 => read_data_o <= x"2020";
when 5747 => read_data_o <= x"1818";
when 5748 => read_data_o <= x"e8e8";
when 5749 => read_data_o <= x"0101";
when 5750 => read_data_o <= x"e8e8";
when 5751 => read_data_o <= x"6464";
when 5752 => read_data_o <= x"0000";
when 5753 => read_data_o <= x"0000";
when 5754 => read_data_o <= x"2020";
when 5755 => read_data_o <= x"0202";
when 5756 => read_data_o <= x"0000";
when 5757 => read_data_o <= x"0000";
when 5758 => read_data_o <= x"0202";
when 5759 => read_data_o <= x"0303";
when 5760 => read_data_o <= x"0101";
when 5761 => read_data_o <= x"0303";
when 5762 => read_data_o <= x"ffff";
when 5763 => read_data_o <= x"a7a7";
when 5764 => read_data_o <= x"0000";
when 5765 => read_data_o <= x"0000";
when 5766 => read_data_o <= x"0000";
when 5767 => read_data_o <= x"0000";
when 5768 => read_data_o <= x"0000";
when 5769 => read_data_o <= x"0000";
when 5770 => read_data_o <= x"0000";
when 5771 => read_data_o <= x"0000";
when 5772 => read_data_o <= x"0000";
when 5773 => read_data_o <= x"0000";
when 5774 => read_data_o <= x"0000";
when 5775 => read_data_o <= x"0000";
when 5776 => read_data_o <= x"0000";
when 5777 => read_data_o <= x"0000";
when 5778 => read_data_o <= x"0000";
when 5779 => read_data_o <= x"0000";
when 5780 => read_data_o <= x"0000";
when 5781 => read_data_o <= x"0000";
when 5782 => read_data_o <= x"0000";
when 5783 => read_data_o <= x"0000";
when 5784 => read_data_o <= x"0000";
when 5785 => read_data_o <= x"0000";
when 5786 => read_data_o <= x"0000";
when 5787 => read_data_o <= x"0000";
when 5788 => read_data_o <= x"0000";
when 5789 => read_data_o <= x"0000";
when 5790 => read_data_o <= x"0000";
when 5791 => read_data_o <= x"0000";
when 5792 => read_data_o <= x"0000";
when 5793 => read_data_o <= x"0000";
when 5794 => read_data_o <= x"0000";
when 5795 => read_data_o <= x"0000";
when 5796 => read_data_o <= x"0000";
when 5797 => read_data_o <= x"0000";
when 5798 => read_data_o <= x"0000";
when 5799 => read_data_o <= x"0000";
when 5800 => read_data_o <= x"0000";
when 5801 => read_data_o <= x"0000";
when 5802 => read_data_o <= x"0000";
when 5803 => read_data_o <= x"0000";
when 5804 => read_data_o <= x"0000";
when 5805 => read_data_o <= x"0000";
when 5806 => read_data_o <= x"0000";
when 5807 => read_data_o <= x"0000";
when 5808 => read_data_o <= x"0000";
when 5809 => read_data_o <= x"0000";
when 5810 => read_data_o <= x"0000";
when 5811 => read_data_o <= x"0000";
when 5812 => read_data_o <= x"d770";
when 5813 => read_data_o <= x"041a";
when 5814 => read_data_o <= x"0000";
when 5815 => read_data_o <= x"0000";
when 5816 => read_data_o <= x"000e";
when 5817 => read_data_o <= x"0000";
when 5818 => read_data_o <= x"0000";
when 5819 => read_data_o <= x"0000";
when 5820 => read_data_o <= x"0000";
when 5821 => read_data_o <= x"0000";
when 5822 => read_data_o <= x"2200";
when 5823 => read_data_o <= x"45d1";
when 5824 => read_data_o <= x"0000";
when 5825 => read_data_o <= x"0000";
when 5826 => read_data_o <= x"0000";
when 5827 => read_data_o <= x"0000";
when 5828 => read_data_o <= x"0000";
when 5829 => read_data_o <= x"0000";
when 5830 => read_data_o <= x"0000";
when 5831 => read_data_o <= x"0000";
when 5832 => read_data_o <= x"0000";
when 5833 => read_data_o <= x"0000";
when 5834 => read_data_o <= x"0000";
when 5835 => read_data_o <= x"0000";
when 5836 => read_data_o <= x"0000";
when 5837 => read_data_o <= x"0000";
when 5838 => read_data_o <= x"0000";
when 5839 => read_data_o <= x"0000";
when 5840 => read_data_o <= x"0000";
when 5841 => read_data_o <= x"0000";
when 5842 => read_data_o <= x"0000";
when 5843 => read_data_o <= x"0000";
when 5844 => read_data_o <= x"0000";
when 5845 => read_data_o <= x"0000";
when 5846 => read_data_o <= x"0000";
when 5847 => read_data_o <= x"0000";
when 5848 => read_data_o <= x"0000";
when 5849 => read_data_o <= x"0000";
when 5850 => read_data_o <= x"0000";
when 5851 => read_data_o <= x"0000";
when 5852 => read_data_o <= x"0000";
when 5853 => read_data_o <= x"0000";
when 5854 => read_data_o <= x"0000";
when 5855 => read_data_o <= x"0000";
when 5856 => read_data_o <= x"0000";
when 5857 => read_data_o <= x"0000";
when 5858 => read_data_o <= x"0000";
when 5859 => read_data_o <= x"0000";
when 5860 => read_data_o <= x"0000";
when 5861 => read_data_o <= x"0000";
when 5862 => read_data_o <= x"0000";
when 5863 => read_data_o <= x"0000";
when 5864 => read_data_o <= x"0000";
when 5865 => read_data_o <= x"0000";
when 5866 => read_data_o <= x"0000";
when 5867 => read_data_o <= x"0000";
when 5868 => read_data_o <= x"0000";
when 5869 => read_data_o <= x"0000";
when 5870 => read_data_o <= x"0000";
when 5871 => read_data_o <= x"0000";
when 5872 => read_data_o <= x"0000";
when 5873 => read_data_o <= x"0000";
when 5874 => read_data_o <= x"0000";
when 5875 => read_data_o <= x"0000";
when 5876 => read_data_o <= x"0000";
when 5877 => read_data_o <= x"0000";
when 5878 => read_data_o <= x"0000";
when 5879 => read_data_o <= x"0000";
when 5880 => read_data_o <= x"0000";
when 5881 => read_data_o <= x"0000";
when 5882 => read_data_o <= x"0000";
when 5883 => read_data_o <= x"0000";
when 5884 => read_data_o <= x"0000";
when 5885 => read_data_o <= x"0000";
when 5886 => read_data_o <= x"0000";
when 5887 => read_data_o <= x"0000";
when 5888 => read_data_o <= x"0000";
when 5889 => read_data_o <= x"0000";
when 5890 => read_data_o <= x"0000";
when 5891 => read_data_o <= x"0000";
when 5892 => read_data_o <= x"d770";
when 5893 => read_data_o <= x"041a";
when 5894 => read_data_o <= x"0000";
when 5895 => read_data_o <= x"0000";
when 5896 => read_data_o <= x"000f";
when 5897 => read_data_o <= x"0000";
when 5898 => read_data_o <= x"0000";
when 5899 => read_data_o <= x"0000";
when 5900 => read_data_o <= x"0000";
when 5901 => read_data_o <= x"0000";
when 5902 => read_data_o <= x"0000";
when 5903 => read_data_o <= x"0000";
when 5904 => read_data_o <= x"0000";
when 5905 => read_data_o <= x"0000";
when 5906 => read_data_o <= x"0000";
when 5907 => read_data_o <= x"0000";
when 5908 => read_data_o <= x"0000";
when 5909 => read_data_o <= x"0000";
when 5910 => read_data_o <= x"0000";
when 5911 => read_data_o <= x"0000";
when 5912 => read_data_o <= x"0000";
when 5913 => read_data_o <= x"0000";
when 5914 => read_data_o <= x"0000";
when 5915 => read_data_o <= x"0000";
when 5916 => read_data_o <= x"0000";
when 5917 => read_data_o <= x"0000";
when 5918 => read_data_o <= x"0000";
when 5919 => read_data_o <= x"0000";
when 5920 => read_data_o <= x"0000";
when 5921 => read_data_o <= x"0000";
when 5922 => read_data_o <= x"0000";
when 5923 => read_data_o <= x"0000";
when 5924 => read_data_o <= x"0000";
when 5925 => read_data_o <= x"0000";
when 5926 => read_data_o <= x"0000";
when 5927 => read_data_o <= x"0000";
when 5928 => read_data_o <= x"0000";
when 5929 => read_data_o <= x"0000";
when 5930 => read_data_o <= x"0000";
when 5931 => read_data_o <= x"0000";
when 5932 => read_data_o <= x"0000";
when 5933 => read_data_o <= x"0000";
when 5934 => read_data_o <= x"0000";
when 5935 => read_data_o <= x"0000";
when 5936 => read_data_o <= x"0000";
when 5937 => read_data_o <= x"0000";
when 5938 => read_data_o <= x"0000";
when 5939 => read_data_o <= x"0000";
when 5940 => read_data_o <= x"0000";
when 5941 => read_data_o <= x"0000";
when 5942 => read_data_o <= x"0000";
when 5943 => read_data_o <= x"0000";
when 5944 => read_data_o <= x"0000";
when 5945 => read_data_o <= x"0000";
when 5946 => read_data_o <= x"0000";
when 5947 => read_data_o <= x"0000";
when 5948 => read_data_o <= x"0000";
when 5949 => read_data_o <= x"0000";
when 5950 => read_data_o <= x"0000";
when 5951 => read_data_o <= x"0000";
when 5952 => read_data_o <= x"0000";
when 5953 => read_data_o <= x"0000";
when 5954 => read_data_o <= x"0000";
when 5955 => read_data_o <= x"0000";
when 5956 => read_data_o <= x"0000";
when 5957 => read_data_o <= x"0000";
when 5958 => read_data_o <= x"0000";
when 5959 => read_data_o <= x"0000";
when 5960 => read_data_o <= x"0000";
when 5961 => read_data_o <= x"0000";
when 5962 => read_data_o <= x"0000";
when 5963 => read_data_o <= x"0000";
when 5964 => read_data_o <= x"0000";
when 5965 => read_data_o <= x"0000";
when 5966 => read_data_o <= x"0000";
when 5967 => read_data_o <= x"0000";
when 5968 => read_data_o <= x"0000";
when 5969 => read_data_o <= x"0000";
when 5970 => read_data_o <= x"0000";
when 5971 => read_data_o <= x"0000";
when 5972 => read_data_o <= x"d770";
when 5973 => read_data_o <= x"041a";
when 5974 => read_data_o <= x"0000";
when 5975 => read_data_o <= x"0000";
when 5976 => read_data_o <= x"0010";
when 5977 => read_data_o <= x"0000";
when 5978 => read_data_o <= x"0000";
when 5979 => read_data_o <= x"0000";
when 5980 => read_data_o <= x"0000";
when 5981 => read_data_o <= x"0000";
when 5982 => read_data_o <= x"0000";
when 5983 => read_data_o <= x"0079";
when 5984 => read_data_o <= x"0000";
when 5985 => read_data_o <= x"0000";
when 5986 => read_data_o <= x"0000";
when 5987 => read_data_o <= x"0000";
when 5988 => read_data_o <= x"0000";
when 5989 => read_data_o <= x"0000";
when 5990 => read_data_o <= x"0000";
when 5991 => read_data_o <= x"0000";
when 5992 => read_data_o <= x"0000";
when 5993 => read_data_o <= x"0000";
when 5994 => read_data_o <= x"0000";
when 5995 => read_data_o <= x"0000";
when 5996 => read_data_o <= x"0000";
when 5997 => read_data_o <= x"0000";
when 5998 => read_data_o <= x"0000";
when 5999 => read_data_o <= x"0000";
when 6000 => read_data_o <= x"0000";
when 6001 => read_data_o <= x"0000";
when 6002 => read_data_o <= x"0000";
when 6003 => read_data_o <= x"0000";
when 6004 => read_data_o <= x"0000";
when 6005 => read_data_o <= x"0000";
when 6006 => read_data_o <= x"0000";
when 6007 => read_data_o <= x"0000";
when 6008 => read_data_o <= x"0000";
when 6009 => read_data_o <= x"0000";
when 6010 => read_data_o <= x"0000";
when 6011 => read_data_o <= x"0000";
when 6012 => read_data_o <= x"0000";
when 6013 => read_data_o <= x"0000";
when 6014 => read_data_o <= x"0000";
when 6015 => read_data_o <= x"0000";
when 6016 => read_data_o <= x"0000";
when 6017 => read_data_o <= x"0000";
when 6018 => read_data_o <= x"0000";
when 6019 => read_data_o <= x"0000";
when 6020 => read_data_o <= x"0000";
when 6021 => read_data_o <= x"0000";
when 6022 => read_data_o <= x"0000";
when 6023 => read_data_o <= x"0000";
when 6024 => read_data_o <= x"0000";
when 6025 => read_data_o <= x"0000";
when 6026 => read_data_o <= x"0000";
when 6027 => read_data_o <= x"0000";
when 6028 => read_data_o <= x"0000";
when 6029 => read_data_o <= x"0000";
when 6030 => read_data_o <= x"0000";
when 6031 => read_data_o <= x"0000";
when 6032 => read_data_o <= x"0000";
when 6033 => read_data_o <= x"0000";
when 6034 => read_data_o <= x"0000";
when 6035 => read_data_o <= x"0000";
when 6036 => read_data_o <= x"0000";
when 6037 => read_data_o <= x"0000";
when 6038 => read_data_o <= x"0000";
when 6039 => read_data_o <= x"0000";
when 6040 => read_data_o <= x"0000";
when 6041 => read_data_o <= x"0000";
when 6042 => read_data_o <= x"0000";
when 6043 => read_data_o <= x"0000";
when 6044 => read_data_o <= x"0000";
when 6045 => read_data_o <= x"0000";
when 6046 => read_data_o <= x"0000";
when 6047 => read_data_o <= x"0000";
when 6048 => read_data_o <= x"0000";
when 6049 => read_data_o <= x"0000";
when 6050 => read_data_o <= x"0000";
when 6051 => read_data_o <= x"0000";
when 6052 => read_data_o <= x"d770";
when 6053 => read_data_o <= x"041a";
when 6054 => read_data_o <= x"0000";
when 6055 => read_data_o <= x"0000";
when 6056 => read_data_o <= x"0011";
when 6057 => read_data_o <= x"0000";
when 6058 => read_data_o <= x"0000";
when 6059 => read_data_o <= x"0000";
when 6060 => read_data_o <= x"0000";
when 6061 => read_data_o <= x"0000";
when 6062 => read_data_o <= x"0000";
when 6063 => read_data_o <= x"0000";
when 6064 => read_data_o <= x"0000";
when 6065 => read_data_o <= x"0000";
when 6066 => read_data_o <= x"0000";
when 6067 => read_data_o <= x"0000";
when 6068 => read_data_o <= x"0000";
when 6069 => read_data_o <= x"0000";
when 6070 => read_data_o <= x"0000";
when 6071 => read_data_o <= x"0000";
when 6072 => read_data_o <= x"0000";
when 6073 => read_data_o <= x"0000";
when 6074 => read_data_o <= x"0000";
when 6075 => read_data_o <= x"0000";
when 6076 => read_data_o <= x"0000";
when 6077 => read_data_o <= x"0000";
when 6078 => read_data_o <= x"0000";
when 6079 => read_data_o <= x"0000";
when 6080 => read_data_o <= x"0000";
when 6081 => read_data_o <= x"0000";
when 6082 => read_data_o <= x"0000";
when 6083 => read_data_o <= x"0000";
when 6084 => read_data_o <= x"0000";
when 6085 => read_data_o <= x"0000";
when 6086 => read_data_o <= x"0000";
when 6087 => read_data_o <= x"0000";
when 6088 => read_data_o <= x"0000";
when 6089 => read_data_o <= x"0000";
when 6090 => read_data_o <= x"0000";
when 6091 => read_data_o <= x"0000";
when 6092 => read_data_o <= x"0000";
when 6093 => read_data_o <= x"0000";
when 6094 => read_data_o <= x"0000";
when 6095 => read_data_o <= x"0000";
when 6096 => read_data_o <= x"0000";
when 6097 => read_data_o <= x"0000";
when 6098 => read_data_o <= x"0000";
when 6099 => read_data_o <= x"0000";
when 6100 => read_data_o <= x"0000";
when 6101 => read_data_o <= x"0000";
when 6102 => read_data_o <= x"0000";
when 6103 => read_data_o <= x"0000";
when 6104 => read_data_o <= x"0000";
when 6105 => read_data_o <= x"0000";
when 6106 => read_data_o <= x"0000";
when 6107 => read_data_o <= x"0000";
when 6108 => read_data_o <= x"0000";
when 6109 => read_data_o <= x"0000";
when 6110 => read_data_o <= x"0000";
when 6111 => read_data_o <= x"0000";
when 6112 => read_data_o <= x"0000";
when 6113 => read_data_o <= x"0000";
when 6114 => read_data_o <= x"0000";
when 6115 => read_data_o <= x"0000";
when 6116 => read_data_o <= x"0000";
when 6117 => read_data_o <= x"0000";
when 6118 => read_data_o <= x"0000";
when 6119 => read_data_o <= x"0000";
when 6120 => read_data_o <= x"0000";
when 6121 => read_data_o <= x"0000";
when 6122 => read_data_o <= x"0000";
when 6123 => read_data_o <= x"0000";
when 6124 => read_data_o <= x"0000";
when 6125 => read_data_o <= x"0000";
when 6126 => read_data_o <= x"0000";
when 6127 => read_data_o <= x"0000";
when 6128 => read_data_o <= x"0000";
when 6129 => read_data_o <= x"0000";
when 6130 => read_data_o <= x"0000";
when 6131 => read_data_o <= x"0000";
when 6132 => read_data_o <= x"d770";
when 6133 => read_data_o <= x"041a";
when 6134 => read_data_o <= x"0000";
when 6135 => read_data_o <= x"0000";
when 6136 => read_data_o <= x"0012";
when 6137 => read_data_o <= x"0000";
when 6138 => read_data_o <= x"0000";
when 6139 => read_data_o <= x"0000";
when 6140 => read_data_o <= x"0000";
when 6141 => read_data_o <= x"0000";
when 6142 => read_data_o <= x"0000";
when 6143 => read_data_o <= x"0000";
when 6144 => read_data_o <= x"0000";
when 6145 => read_data_o <= x"0000";
when 6146 => read_data_o <= x"0000";
when 6147 => read_data_o <= x"0000";
when 6148 => read_data_o <= x"0000";
when 6149 => read_data_o <= x"0000";
when 6150 => read_data_o <= x"0000";
when 6151 => read_data_o <= x"0000";
when 6152 => read_data_o <= x"0000";
when 6153 => read_data_o <= x"0000";
when 6154 => read_data_o <= x"0000";
when 6155 => read_data_o <= x"0000";
when 6156 => read_data_o <= x"0000";
when 6157 => read_data_o <= x"0000";
when 6158 => read_data_o <= x"0000";
when 6159 => read_data_o <= x"0000";
when 6160 => read_data_o <= x"0000";
when 6161 => read_data_o <= x"0000";
when 6162 => read_data_o <= x"0000";
when 6163 => read_data_o <= x"0000";
when 6164 => read_data_o <= x"0000";
when 6165 => read_data_o <= x"0000";
when 6166 => read_data_o <= x"0000";
when 6167 => read_data_o <= x"0000";
when 6168 => read_data_o <= x"0000";
when 6169 => read_data_o <= x"0000";
when 6170 => read_data_o <= x"0000";
when 6171 => read_data_o <= x"0000";
when 6172 => read_data_o <= x"0000";
when 6173 => read_data_o <= x"0000";
when 6174 => read_data_o <= x"0000";
when 6175 => read_data_o <= x"0000";
when 6176 => read_data_o <= x"0000";
when 6177 => read_data_o <= x"0000";
when 6178 => read_data_o <= x"0000";
when 6179 => read_data_o <= x"0000";
when 6180 => read_data_o <= x"0000";
when 6181 => read_data_o <= x"0000";
when 6182 => read_data_o <= x"0000";
when 6183 => read_data_o <= x"0000";
when 6184 => read_data_o <= x"0000";
when 6185 => read_data_o <= x"0000";
when 6186 => read_data_o <= x"0000";
when 6187 => read_data_o <= x"0000";
when 6188 => read_data_o <= x"0000";
when 6189 => read_data_o <= x"0000";
when 6190 => read_data_o <= x"0000";
when 6191 => read_data_o <= x"0000";
when 6192 => read_data_o <= x"0000";
when 6193 => read_data_o <= x"0000";
when 6194 => read_data_o <= x"0000";
when 6195 => read_data_o <= x"0000";
when 6196 => read_data_o <= x"0000";
when 6197 => read_data_o <= x"0000";
when 6198 => read_data_o <= x"0000";
when 6199 => read_data_o <= x"0000";
when 6200 => read_data_o <= x"0000";
when 6201 => read_data_o <= x"0000";
when 6202 => read_data_o <= x"0000";
when 6203 => read_data_o <= x"0000";
when 6204 => read_data_o <= x"0000";
when 6205 => read_data_o <= x"0000";
when 6206 => read_data_o <= x"0000";
when 6207 => read_data_o <= x"0000";
when 6208 => read_data_o <= x"0000";
when 6209 => read_data_o <= x"0000";
when 6210 => read_data_o <= x"0000";
when 6211 => read_data_o <= x"0000";
when 6212 => read_data_o <= x"d770";
when 6213 => read_data_o <= x"041a";
when 6214 => read_data_o <= x"0000";
when 6215 => read_data_o <= x"0000";
when 6216 => read_data_o <= x"0013";
when 6217 => read_data_o <= x"0000";
when 6218 => read_data_o <= x"0000";
when 6219 => read_data_o <= x"0000";
when 6220 => read_data_o <= x"0000";
when 6221 => read_data_o <= x"0000";
when 6222 => read_data_o <= x"0000";
when 6223 => read_data_o <= x"0000";
when 6224 => read_data_o <= x"0000";
when 6225 => read_data_o <= x"0000";
when 6226 => read_data_o <= x"0000";
when 6227 => read_data_o <= x"0000";
when 6228 => read_data_o <= x"0000";
when 6229 => read_data_o <= x"0000";
when 6230 => read_data_o <= x"0000";
when 6231 => read_data_o <= x"0000";
when 6232 => read_data_o <= x"0000";
when 6233 => read_data_o <= x"0000";
when 6234 => read_data_o <= x"0000";
when 6235 => read_data_o <= x"0000";
when 6236 => read_data_o <= x"0000";
when 6237 => read_data_o <= x"0000";
when 6238 => read_data_o <= x"0000";
when 6239 => read_data_o <= x"0000";
when 6240 => read_data_o <= x"0000";
when 6241 => read_data_o <= x"0000";
when 6242 => read_data_o <= x"0000";
when 6243 => read_data_o <= x"0000";
when 6244 => read_data_o <= x"0000";
when 6245 => read_data_o <= x"0000";
when 6246 => read_data_o <= x"0000";
when 6247 => read_data_o <= x"0000";
when 6248 => read_data_o <= x"0000";
when 6249 => read_data_o <= x"0000";
when 6250 => read_data_o <= x"0000";
when 6251 => read_data_o <= x"0000";
when 6252 => read_data_o <= x"0000";
when 6253 => read_data_o <= x"0000";
when 6254 => read_data_o <= x"0000";
when 6255 => read_data_o <= x"0000";
when 6256 => read_data_o <= x"0000";
when 6257 => read_data_o <= x"0000";
when 6258 => read_data_o <= x"0000";
when 6259 => read_data_o <= x"0000";
when 6260 => read_data_o <= x"0000";
when 6261 => read_data_o <= x"0000";
when 6262 => read_data_o <= x"0000";
when 6263 => read_data_o <= x"0000";
when 6264 => read_data_o <= x"0000";
when 6265 => read_data_o <= x"0000";
when 6266 => read_data_o <= x"0000";
when 6267 => read_data_o <= x"0000";
when 6268 => read_data_o <= x"0000";
when 6269 => read_data_o <= x"0000";
when 6270 => read_data_o <= x"0000";
when 6271 => read_data_o <= x"0000";
when 6272 => read_data_o <= x"0000";
when 6273 => read_data_o <= x"0000";
when 6274 => read_data_o <= x"0000";
when 6275 => read_data_o <= x"0000";
when 6276 => read_data_o <= x"0000";
when 6277 => read_data_o <= x"0000";
when 6278 => read_data_o <= x"0000";
when 6279 => read_data_o <= x"0000";
when 6280 => read_data_o <= x"0000";
when 6281 => read_data_o <= x"0000";
when 6282 => read_data_o <= x"0000";
when 6283 => read_data_o <= x"0000";
when 6284 => read_data_o <= x"0000";
when 6285 => read_data_o <= x"0000";
when 6286 => read_data_o <= x"0000";
when 6287 => read_data_o <= x"0000";
when 6288 => read_data_o <= x"0000";
when 6289 => read_data_o <= x"0000";
when 6290 => read_data_o <= x"0000";
when 6291 => read_data_o <= x"0000";
when 6292 => read_data_o <= x"d770";
when 6293 => read_data_o <= x"041a";
when 6294 => read_data_o <= x"0000";
when 6295 => read_data_o <= x"0000";
when 6296 => read_data_o <= x"0014";
when 6297 => read_data_o <= x"0000";
when 6298 => read_data_o <= x"0000";
when 6299 => read_data_o <= x"0000";
when 6300 => read_data_o <= x"0000";
when 6301 => read_data_o <= x"0000";
when 6302 => read_data_o <= x"0000";
when 6303 => read_data_o <= x"0000";
when 6304 => read_data_o <= x"0000";
when 6305 => read_data_o <= x"0000";
when 6306 => read_data_o <= x"0000";
when 6307 => read_data_o <= x"0000";
when 6308 => read_data_o <= x"0000";
when 6309 => read_data_o <= x"0000";
when 6310 => read_data_o <= x"0000";
when 6311 => read_data_o <= x"0000";
when 6312 => read_data_o <= x"0000";
when 6313 => read_data_o <= x"0000";
when 6314 => read_data_o <= x"0000";
when 6315 => read_data_o <= x"0000";
when 6316 => read_data_o <= x"0000";
when 6317 => read_data_o <= x"0000";
when 6318 => read_data_o <= x"0000";
when 6319 => read_data_o <= x"0000";
when 6320 => read_data_o <= x"0000";
when 6321 => read_data_o <= x"0000";
when 6322 => read_data_o <= x"0000";
when 6323 => read_data_o <= x"0000";
when 6324 => read_data_o <= x"0000";
when 6325 => read_data_o <= x"0000";
when 6326 => read_data_o <= x"0000";
when 6327 => read_data_o <= x"0000";
when 6328 => read_data_o <= x"0000";
when 6329 => read_data_o <= x"0000";
when 6330 => read_data_o <= x"0000";
when 6331 => read_data_o <= x"0000";
when 6332 => read_data_o <= x"0000";
when 6333 => read_data_o <= x"0000";
when 6334 => read_data_o <= x"0000";
when 6335 => read_data_o <= x"0000";
when 6336 => read_data_o <= x"0000";
when 6337 => read_data_o <= x"0000";
when 6338 => read_data_o <= x"0000";
when 6339 => read_data_o <= x"0000";
when 6340 => read_data_o <= x"0000";
when 6341 => read_data_o <= x"0000";
when 6342 => read_data_o <= x"0000";
when 6343 => read_data_o <= x"0000";
when 6344 => read_data_o <= x"0000";
when 6345 => read_data_o <= x"0000";
when 6346 => read_data_o <= x"0000";
when 6347 => read_data_o <= x"0000";
when 6348 => read_data_o <= x"0000";
when 6349 => read_data_o <= x"0000";
when 6350 => read_data_o <= x"0000";
when 6351 => read_data_o <= x"0000";
when 6352 => read_data_o <= x"0000";
when 6353 => read_data_o <= x"0000";
when 6354 => read_data_o <= x"0000";
when 6355 => read_data_o <= x"0000";
when 6356 => read_data_o <= x"0000";
when 6357 => read_data_o <= x"0000";
when 6358 => read_data_o <= x"0000";
when 6359 => read_data_o <= x"0000";
when 6360 => read_data_o <= x"0000";
when 6361 => read_data_o <= x"0000";
when 6362 => read_data_o <= x"0000";
when 6363 => read_data_o <= x"0000";
when 6364 => read_data_o <= x"0000";
when 6365 => read_data_o <= x"0000";
when 6366 => read_data_o <= x"0000";
when 6367 => read_data_o <= x"0000";
when 6368 => read_data_o <= x"0000";
when 6369 => read_data_o <= x"0000";
when 6370 => read_data_o <= x"0000";
when 6371 => read_data_o <= x"0000";
when 6372 => read_data_o <= x"d770";
when 6373 => read_data_o <= x"041a";
when 6374 => read_data_o <= x"0000";
when 6375 => read_data_o <= x"0000";
when 6376 => read_data_o <= x"0015";
when 6377 => read_data_o <= x"0000";
when 6378 => read_data_o <= x"0000";
when 6379 => read_data_o <= x"0000";
when 6380 => read_data_o <= x"0000";
when 6381 => read_data_o <= x"0000";
when 6382 => read_data_o <= x"0000";
when 6383 => read_data_o <= x"0000";
when 6384 => read_data_o <= x"0000";
when 6385 => read_data_o <= x"0000";
when 6386 => read_data_o <= x"0000";
when 6387 => read_data_o <= x"0000";
when 6388 => read_data_o <= x"0000";
when 6389 => read_data_o <= x"0000";
when 6390 => read_data_o <= x"0000";
when 6391 => read_data_o <= x"0000";
when 6392 => read_data_o <= x"0000";
when 6393 => read_data_o <= x"0000";
when 6394 => read_data_o <= x"0000";
when 6395 => read_data_o <= x"0000";
when 6396 => read_data_o <= x"0000";
when 6397 => read_data_o <= x"0000";
when 6398 => read_data_o <= x"0000";
when 6399 => read_data_o <= x"0000";
when 6400 => read_data_o <= x"0000";
when 6401 => read_data_o <= x"0000";
when 6402 => read_data_o <= x"0000";
when 6403 => read_data_o <= x"0000";
when 6404 => read_data_o <= x"0000";
when 6405 => read_data_o <= x"0000";
when 6406 => read_data_o <= x"0000";
when 6407 => read_data_o <= x"0000";
when 6408 => read_data_o <= x"0000";
when 6409 => read_data_o <= x"0000";
when 6410 => read_data_o <= x"0000";
when 6411 => read_data_o <= x"0000";
when 6412 => read_data_o <= x"0000";
when 6413 => read_data_o <= x"0000";
when 6414 => read_data_o <= x"0000";
when 6415 => read_data_o <= x"0000";
when 6416 => read_data_o <= x"0000";
when 6417 => read_data_o <= x"0000";
when 6418 => read_data_o <= x"0000";
when 6419 => read_data_o <= x"0000";
when 6420 => read_data_o <= x"0000";
when 6421 => read_data_o <= x"0000";
when 6422 => read_data_o <= x"0000";
when 6423 => read_data_o <= x"0000";
when 6424 => read_data_o <= x"0000";
when 6425 => read_data_o <= x"0000";
when 6426 => read_data_o <= x"0000";
when 6427 => read_data_o <= x"0000";
when 6428 => read_data_o <= x"0000";
when 6429 => read_data_o <= x"0000";
when 6430 => read_data_o <= x"0000";
when 6431 => read_data_o <= x"0000";
when 6432 => read_data_o <= x"0000";
when 6433 => read_data_o <= x"0000";
when 6434 => read_data_o <= x"0000";
when 6435 => read_data_o <= x"0000";
when 6436 => read_data_o <= x"0000";
when 6437 => read_data_o <= x"0000";
when 6438 => read_data_o <= x"0000";
when 6439 => read_data_o <= x"0000";
when 6440 => read_data_o <= x"0000";
when 6441 => read_data_o <= x"0000";
when 6442 => read_data_o <= x"0000";
when 6443 => read_data_o <= x"0000";
when 6444 => read_data_o <= x"0000";
when 6445 => read_data_o <= x"0000";
when 6446 => read_data_o <= x"0000";
when 6447 => read_data_o <= x"0000";
when 6448 => read_data_o <= x"0000";
when 6449 => read_data_o <= x"0000";
when 6450 => read_data_o <= x"0032";
when 6451 => read_data_o <= x"2e30";
when 6452 => read_data_o <= x"d770";
when 6453 => read_data_o <= x"041a";
when 6454 => read_data_o <= x"0000";
when 6455 => read_data_o <= x"0000";
when 6456 => read_data_o <= x"0016";
when 6457 => read_data_o <= x"0000";
when 6458 => read_data_o <= x"0000";
when 6459 => read_data_o <= x"0000";
when 6460 => read_data_o <= x"0000";
when 6461 => read_data_o <= x"0000";
when 6462 => read_data_o <= x"0000";
when 6463 => read_data_o <= x"0000";
when 6464 => read_data_o <= x"0000";
when 6465 => read_data_o <= x"0000";
when 6466 => read_data_o <= x"0000";
when 6467 => read_data_o <= x"0000";
when 6468 => read_data_o <= x"0000";
when 6469 => read_data_o <= x"0000";
when 6470 => read_data_o <= x"0000";
when 6471 => read_data_o <= x"0000";
when 6472 => read_data_o <= x"0000";
when 6473 => read_data_o <= x"0000";
when 6474 => read_data_o <= x"0000";
when 6475 => read_data_o <= x"0000";
when 6476 => read_data_o <= x"0000";
when 6477 => read_data_o <= x"0000";
when 6478 => read_data_o <= x"0000";
when 6479 => read_data_o <= x"0000";
when 6480 => read_data_o <= x"0000";
when 6481 => read_data_o <= x"0000";
when 6482 => read_data_o <= x"0000";
when 6483 => read_data_o <= x"0000";
when 6484 => read_data_o <= x"0000";
when 6485 => read_data_o <= x"0000";
when 6486 => read_data_o <= x"0000";
when 6487 => read_data_o <= x"0000";
when 6488 => read_data_o <= x"0000";
when 6489 => read_data_o <= x"0000";
when 6490 => read_data_o <= x"0000";
when 6491 => read_data_o <= x"0000";
when 6492 => read_data_o <= x"0000";
when 6493 => read_data_o <= x"0000";
when 6494 => read_data_o <= x"0000";
when 6495 => read_data_o <= x"0000";
when 6496 => read_data_o <= x"0000";
when 6497 => read_data_o <= x"0000";
when 6498 => read_data_o <= x"0000";
when 6499 => read_data_o <= x"0000";
when 6500 => read_data_o <= x"0000";
when 6501 => read_data_o <= x"0000";
when 6502 => read_data_o <= x"0000";
when 6503 => read_data_o <= x"0000";
when 6504 => read_data_o <= x"0000";
when 6505 => read_data_o <= x"0000";
when 6506 => read_data_o <= x"0000";
when 6507 => read_data_o <= x"0000";
when 6508 => read_data_o <= x"0000";
when 6509 => read_data_o <= x"0000";
when 6510 => read_data_o <= x"0000";
when 6511 => read_data_o <= x"0000";
when 6512 => read_data_o <= x"0000";
when 6513 => read_data_o <= x"0000";
when 6514 => read_data_o <= x"0000";
when 6515 => read_data_o <= x"0000";
when 6516 => read_data_o <= x"0000";
when 6517 => read_data_o <= x"0000";
when 6518 => read_data_o <= x"0000";
when 6519 => read_data_o <= x"0000";
when 6520 => read_data_o <= x"0000";
when 6521 => read_data_o <= x"0000";
when 6522 => read_data_o <= x"0000";
when 6523 => read_data_o <= x"0000";
when 6524 => read_data_o <= x"0000";
when 6525 => read_data_o <= x"0000";
when 6526 => read_data_o <= x"0000";
when 6527 => read_data_o <= x"0000";
when 6528 => read_data_o <= x"0000";
when 6529 => read_data_o <= x"0000";
when 6530 => read_data_o <= x"0000";
when 6531 => read_data_o <= x"0000";
when 6532 => read_data_o <= x"d770";
when 6533 => read_data_o <= x"041a";
when 6534 => read_data_o <= x"0000";
when 6535 => read_data_o <= x"0000";
when 6536 => read_data_o <= x"0017";
when 6537 => read_data_o <= x"0000";
when 6538 => read_data_o <= x"0000";
when 6539 => read_data_o <= x"0000";
when 6540 => read_data_o <= x"0000";
when 6541 => read_data_o <= x"0000";
when 6542 => read_data_o <= x"6500";
when 6543 => read_data_o <= x"0000";
when 6544 => read_data_o <= x"0000";
when 6545 => read_data_o <= x"0000";
when 6546 => read_data_o <= x"0000";
when 6547 => read_data_o <= x"0000";
when 6548 => read_data_o <= x"0000";
when 6549 => read_data_o <= x"0000";
when 6550 => read_data_o <= x"0000";
when 6551 => read_data_o <= x"0000";
when 6552 => read_data_o <= x"0000";
when 6553 => read_data_o <= x"0000";
when 6554 => read_data_o <= x"0000";
when 6555 => read_data_o <= x"0000";
when 6556 => read_data_o <= x"0000";
when 6557 => read_data_o <= x"0000";
when 6558 => read_data_o <= x"0000";
when 6559 => read_data_o <= x"0000";
when 6560 => read_data_o <= x"0000";
when 6561 => read_data_o <= x"0000";
when 6562 => read_data_o <= x"0000";
when 6563 => read_data_o <= x"0000";
when 6564 => read_data_o <= x"0000";
when 6565 => read_data_o <= x"0000";
when 6566 => read_data_o <= x"0000";
when 6567 => read_data_o <= x"0000";
when 6568 => read_data_o <= x"0000";
when 6569 => read_data_o <= x"0000";
when 6570 => read_data_o <= x"0000";
when 6571 => read_data_o <= x"0000";
when 6572 => read_data_o <= x"0000";
when 6573 => read_data_o <= x"0000";
when 6574 => read_data_o <= x"0000";
when 6575 => read_data_o <= x"0000";
when 6576 => read_data_o <= x"0000";
when 6577 => read_data_o <= x"0000";
when 6578 => read_data_o <= x"0000";
when 6579 => read_data_o <= x"0000";
when 6580 => read_data_o <= x"0000";
when 6581 => read_data_o <= x"0000";
when 6582 => read_data_o <= x"0000";
when 6583 => read_data_o <= x"0000";
when 6584 => read_data_o <= x"0000";
when 6585 => read_data_o <= x"0000";
when 6586 => read_data_o <= x"0000";
when 6587 => read_data_o <= x"0000";
when 6588 => read_data_o <= x"0000";
when 6589 => read_data_o <= x"0000";
when 6590 => read_data_o <= x"0000";
when 6591 => read_data_o <= x"0000";
when 6592 => read_data_o <= x"0000";
when 6593 => read_data_o <= x"0000";
when 6594 => read_data_o <= x"0000";
when 6595 => read_data_o <= x"0000";
when 6596 => read_data_o <= x"0000";
when 6597 => read_data_o <= x"0000";
when 6598 => read_data_o <= x"0000";
when 6599 => read_data_o <= x"0000";
when 6600 => read_data_o <= x"0000";
when 6601 => read_data_o <= x"0000";
when 6602 => read_data_o <= x"0000";
when 6603 => read_data_o <= x"0000";
when 6604 => read_data_o <= x"0000";
when 6605 => read_data_o <= x"0000";
when 6606 => read_data_o <= x"0000";
when 6607 => read_data_o <= x"0000";
when 6608 => read_data_o <= x"0000";
when 6609 => read_data_o <= x"0000";
when 6610 => read_data_o <= x"0000";
when 6611 => read_data_o <= x"0000";
when 6612 => read_data_o <= x"d770";
when 6613 => read_data_o <= x"041a";
when 6614 => read_data_o <= x"0000";
when 6615 => read_data_o <= x"0000";
when 6616 => read_data_o <= x"0018";
when 6617 => read_data_o <= x"0000";
when 6618 => read_data_o <= x"0000";
when 6619 => read_data_o <= x"0000";
when 6620 => read_data_o <= x"0000";
when 6621 => read_data_o <= x"0000";
when 6622 => read_data_o <= x"7f00";
when 6623 => read_data_o <= x"0000";
when 6624 => read_data_o <= x"0000";
when 6625 => read_data_o <= x"0000";
when 6626 => read_data_o <= x"0000";
when 6627 => read_data_o <= x"0000";
when 6628 => read_data_o <= x"0000";
when 6629 => read_data_o <= x"0000";
when 6630 => read_data_o <= x"0000";
when 6631 => read_data_o <= x"0000";
when 6632 => read_data_o <= x"0000";
when 6633 => read_data_o <= x"0000";
when 6634 => read_data_o <= x"0000";
when 6635 => read_data_o <= x"0000";
when 6636 => read_data_o <= x"0000";
when 6637 => read_data_o <= x"0000";
when 6638 => read_data_o <= x"0000";
when 6639 => read_data_o <= x"0000";
when 6640 => read_data_o <= x"0000";
when 6641 => read_data_o <= x"0000";
when 6642 => read_data_o <= x"0000";
when 6643 => read_data_o <= x"0000";
when 6644 => read_data_o <= x"0000";
when 6645 => read_data_o <= x"0000";
when 6646 => read_data_o <= x"0000";
when 6647 => read_data_o <= x"0000";
when 6648 => read_data_o <= x"0000";
when 6649 => read_data_o <= x"0000";
when 6650 => read_data_o <= x"0000";
when 6651 => read_data_o <= x"0000";
when 6652 => read_data_o <= x"0000";
when 6653 => read_data_o <= x"0000";
when 6654 => read_data_o <= x"0000";
when 6655 => read_data_o <= x"0000";
when 6656 => read_data_o <= x"0000";
when 6657 => read_data_o <= x"0000";
when 6658 => read_data_o <= x"0000";
when 6659 => read_data_o <= x"0000";
when 6660 => read_data_o <= x"0000";
when 6661 => read_data_o <= x"0000";
when 6662 => read_data_o <= x"0000";
when 6663 => read_data_o <= x"0000";
when 6664 => read_data_o <= x"0000";
when 6665 => read_data_o <= x"0000";
when 6666 => read_data_o <= x"0000";
when 6667 => read_data_o <= x"0000";
when 6668 => read_data_o <= x"0000";
when 6669 => read_data_o <= x"0000";
when 6670 => read_data_o <= x"0000";
when 6671 => read_data_o <= x"0000";
when 6672 => read_data_o <= x"0000";
when 6673 => read_data_o <= x"0000";
when 6674 => read_data_o <= x"0000";
when 6675 => read_data_o <= x"0000";
when 6676 => read_data_o <= x"0000";
when 6677 => read_data_o <= x"0000";
when 6678 => read_data_o <= x"0000";
when 6679 => read_data_o <= x"0000";
when 6680 => read_data_o <= x"0000";
when 6681 => read_data_o <= x"0000";
when 6682 => read_data_o <= x"0000";
when 6683 => read_data_o <= x"0000";
when 6684 => read_data_o <= x"0000";
when 6685 => read_data_o <= x"0000";
when 6686 => read_data_o <= x"0000";
when 6687 => read_data_o <= x"0000";
when 6688 => read_data_o <= x"0000";
when 6689 => read_data_o <= x"0000";
when 6690 => read_data_o <= x"0000";
when 6691 => read_data_o <= x"0000";
when 6692 => read_data_o <= x"d770";
when 6693 => read_data_o <= x"041a";
when 6694 => read_data_o <= x"0000";
when 6695 => read_data_o <= x"0000";
when 6696 => read_data_o <= x"0019";
when 6697 => read_data_o <= x"0000";
when 6698 => read_data_o <= x"0000";
when 6699 => read_data_o <= x"0000";
when 6700 => read_data_o <= x"0000";
when 6701 => read_data_o <= x"0000";
when 6702 => read_data_o <= x"0000";
when 6703 => read_data_o <= x"0000";
when 6704 => read_data_o <= x"0000";
when 6705 => read_data_o <= x"0000";
when 6706 => read_data_o <= x"0000";
when 6707 => read_data_o <= x"0000";
when 6708 => read_data_o <= x"0000";
when 6709 => read_data_o <= x"0000";
when 6710 => read_data_o <= x"0000";
when 6711 => read_data_o <= x"0000";
when 6712 => read_data_o <= x"0000";
when 6713 => read_data_o <= x"0000";
when 6714 => read_data_o <= x"0000";
when 6715 => read_data_o <= x"0000";
when 6716 => read_data_o <= x"0000";
when 6717 => read_data_o <= x"0000";
when 6718 => read_data_o <= x"0000";
when 6719 => read_data_o <= x"0000";
when 6720 => read_data_o <= x"0000";
when 6721 => read_data_o <= x"0000";
when 6722 => read_data_o <= x"0000";
when 6723 => read_data_o <= x"0000";
when 6724 => read_data_o <= x"0000";
when 6725 => read_data_o <= x"0000";
when 6726 => read_data_o <= x"0000";
when 6727 => read_data_o <= x"0000";
when 6728 => read_data_o <= x"0000";
when 6729 => read_data_o <= x"0000";
when 6730 => read_data_o <= x"0000";
when 6731 => read_data_o <= x"0000";
when 6732 => read_data_o <= x"0000";
when 6733 => read_data_o <= x"0000";
when 6734 => read_data_o <= x"0000";
when 6735 => read_data_o <= x"0000";
when 6736 => read_data_o <= x"0000";
when 6737 => read_data_o <= x"0000";
when 6738 => read_data_o <= x"0000";
when 6739 => read_data_o <= x"0000";
when 6740 => read_data_o <= x"0000";
when 6741 => read_data_o <= x"0000";
when 6742 => read_data_o <= x"0000";
when 6743 => read_data_o <= x"0000";
when 6744 => read_data_o <= x"0000";
when 6745 => read_data_o <= x"0000";
when 6746 => read_data_o <= x"0000";
when 6747 => read_data_o <= x"0000";
when 6748 => read_data_o <= x"0000";
when 6749 => read_data_o <= x"0000";
when 6750 => read_data_o <= x"0000";
when 6751 => read_data_o <= x"0000";
when 6752 => read_data_o <= x"0000";
when 6753 => read_data_o <= x"0000";
when 6754 => read_data_o <= x"0000";
when 6755 => read_data_o <= x"0000";
when 6756 => read_data_o <= x"0000";
when 6757 => read_data_o <= x"0000";
when 6758 => read_data_o <= x"0000";
when 6759 => read_data_o <= x"0000";
when 6760 => read_data_o <= x"0000";
when 6761 => read_data_o <= x"0000";
when 6762 => read_data_o <= x"0000";
when 6763 => read_data_o <= x"0000";
when 6764 => read_data_o <= x"0000";
when 6765 => read_data_o <= x"0000";
when 6766 => read_data_o <= x"0000";
when 6767 => read_data_o <= x"0000";
when 6768 => read_data_o <= x"0000";
when 6769 => read_data_o <= x"0000";
when 6770 => read_data_o <= x"0000";
when 6771 => read_data_o <= x"0000";
when 6772 => read_data_o <= x"d770";
when 6773 => read_data_o <= x"041a";
when 6774 => read_data_o <= x"0000";
when 6775 => read_data_o <= x"0000";
when 6776 => read_data_o <= x"001a";
when 6777 => read_data_o <= x"0000";
when 6778 => read_data_o <= x"0000";
when 6779 => read_data_o <= x"0000";
when 6780 => read_data_o <= x"0000";
when 6781 => read_data_o <= x"0000";
when 6782 => read_data_o <= x"0000";
when 6783 => read_data_o <= x"0000";
when 6784 => read_data_o <= x"0000";
when 6785 => read_data_o <= x"0000";
when 6786 => read_data_o <= x"0000";
when 6787 => read_data_o <= x"0000";
when 6788 => read_data_o <= x"0000";
when 6789 => read_data_o <= x"0000";
when 6790 => read_data_o <= x"0000";
when 6791 => read_data_o <= x"0000";
when 6792 => read_data_o <= x"0000";
when 6793 => read_data_o <= x"0000";
when 6794 => read_data_o <= x"0000";
when 6795 => read_data_o <= x"0000";
when 6796 => read_data_o <= x"0000";
when 6797 => read_data_o <= x"0000";
when 6798 => read_data_o <= x"0000";
when 6799 => read_data_o <= x"0000";
when 6800 => read_data_o <= x"0000";
when 6801 => read_data_o <= x"0000";
when 6802 => read_data_o <= x"0000";
when 6803 => read_data_o <= x"0000";
when 6804 => read_data_o <= x"0000";
when 6805 => read_data_o <= x"0000";
when 6806 => read_data_o <= x"0000";
when 6807 => read_data_o <= x"0000";
when 6808 => read_data_o <= x"0000";
when 6809 => read_data_o <= x"0000";
when 6810 => read_data_o <= x"0000";
when 6811 => read_data_o <= x"0000";
when 6812 => read_data_o <= x"0000";
when 6813 => read_data_o <= x"0000";
when 6814 => read_data_o <= x"0000";
when 6815 => read_data_o <= x"0000";
when 6816 => read_data_o <= x"0000";
when 6817 => read_data_o <= x"0000";
when 6818 => read_data_o <= x"0000";
when 6819 => read_data_o <= x"0000";
when 6820 => read_data_o <= x"0000";
when 6821 => read_data_o <= x"0000";
when 6822 => read_data_o <= x"0000";
when 6823 => read_data_o <= x"0000";
when 6824 => read_data_o <= x"0000";
when 6825 => read_data_o <= x"0000";
when 6826 => read_data_o <= x"0000";
when 6827 => read_data_o <= x"0000";
when 6828 => read_data_o <= x"0000";
when 6829 => read_data_o <= x"0000";
when 6830 => read_data_o <= x"0000";
when 6831 => read_data_o <= x"0000";
when 6832 => read_data_o <= x"0000";
when 6833 => read_data_o <= x"0000";
when 6834 => read_data_o <= x"0000";
when 6835 => read_data_o <= x"0000";
when 6836 => read_data_o <= x"0000";
when 6837 => read_data_o <= x"0000";
when 6838 => read_data_o <= x"0000";
when 6839 => read_data_o <= x"0000";
when 6840 => read_data_o <= x"0000";
when 6841 => read_data_o <= x"0000";
when 6842 => read_data_o <= x"0000";
when 6843 => read_data_o <= x"0000";
when 6844 => read_data_o <= x"0000";
when 6845 => read_data_o <= x"0000";
when 6846 => read_data_o <= x"0000";
when 6847 => read_data_o <= x"0000";
when 6848 => read_data_o <= x"0000";
when 6849 => read_data_o <= x"0000";
when 6850 => read_data_o <= x"0000";
when 6851 => read_data_o <= x"0000";
when 6852 => read_data_o <= x"d770";
when 6853 => read_data_o <= x"041a";
when 6854 => read_data_o <= x"0000";
when 6855 => read_data_o <= x"0000";
when 6856 => read_data_o <= x"001b";
when 6857 => read_data_o <= x"0000";
when 6858 => read_data_o <= x"0000";
when 6859 => read_data_o <= x"0000";
when 6860 => read_data_o <= x"0000";
when 6861 => read_data_o <= x"0000";
when 6862 => read_data_o <= x"0000";
when 6863 => read_data_o <= x"0000";
when 6864 => read_data_o <= x"0000";
when 6865 => read_data_o <= x"0000";
when 6866 => read_data_o <= x"0000";
when 6867 => read_data_o <= x"0000";
when 6868 => read_data_o <= x"0000";
when 6869 => read_data_o <= x"0000";
when 6870 => read_data_o <= x"0000";
when 6871 => read_data_o <= x"0000";
when 6872 => read_data_o <= x"0000";
when 6873 => read_data_o <= x"0000";
when 6874 => read_data_o <= x"0000";
when 6875 => read_data_o <= x"0000";
when 6876 => read_data_o <= x"0000";
when 6877 => read_data_o <= x"0000";
when 6878 => read_data_o <= x"0000";
when 6879 => read_data_o <= x"0000";
when 6880 => read_data_o <= x"0000";
when 6881 => read_data_o <= x"0000";
when 6882 => read_data_o <= x"0000";
when 6883 => read_data_o <= x"0000";
when 6884 => read_data_o <= x"0000";
when 6885 => read_data_o <= x"0000";
when 6886 => read_data_o <= x"0000";
when 6887 => read_data_o <= x"0000";
when 6888 => read_data_o <= x"0000";
when 6889 => read_data_o <= x"0000";
when 6890 => read_data_o <= x"0000";
when 6891 => read_data_o <= x"0000";
when 6892 => read_data_o <= x"0000";
when 6893 => read_data_o <= x"0000";
when 6894 => read_data_o <= x"0000";
when 6895 => read_data_o <= x"0000";
when 6896 => read_data_o <= x"0000";
when 6897 => read_data_o <= x"0000";
when 6898 => read_data_o <= x"0000";
when 6899 => read_data_o <= x"0000";
when 6900 => read_data_o <= x"0000";
when 6901 => read_data_o <= x"0000";
when 6902 => read_data_o <= x"0000";
when 6903 => read_data_o <= x"0000";
when 6904 => read_data_o <= x"0000";
when 6905 => read_data_o <= x"0000";
when 6906 => read_data_o <= x"0000";
when 6907 => read_data_o <= x"0000";
when 6908 => read_data_o <= x"0000";
when 6909 => read_data_o <= x"0000";
when 6910 => read_data_o <= x"0000";
when 6911 => read_data_o <= x"0000";
when 6912 => read_data_o <= x"0000";
when 6913 => read_data_o <= x"0000";
when 6914 => read_data_o <= x"0000";
when 6915 => read_data_o <= x"0000";
when 6916 => read_data_o <= x"0000";
when 6917 => read_data_o <= x"0000";
when 6918 => read_data_o <= x"0000";
when 6919 => read_data_o <= x"0000";
when 6920 => read_data_o <= x"0000";
when 6921 => read_data_o <= x"0000";
when 6922 => read_data_o <= x"0000";
when 6923 => read_data_o <= x"0000";
when 6924 => read_data_o <= x"0000";
when 6925 => read_data_o <= x"0000";
when 6926 => read_data_o <= x"0000";
when 6927 => read_data_o <= x"0000";
when 6928 => read_data_o <= x"0000";
when 6929 => read_data_o <= x"0000";
when 6930 => read_data_o <= x"665f";
when 6931 => read_data_o <= x"6172";
when 6932 => read_data_o <= x"d770";
when 6933 => read_data_o <= x"041a";
when 6934 => read_data_o <= x"0000";
when 6935 => read_data_o <= x"0000";
when 6936 => read_data_o <= x"001c";
when 6937 => read_data_o <= x"0000";
when 6938 => read_data_o <= x"0000";
when 6939 => read_data_o <= x"0000";
when 6940 => read_data_o <= x"0000";
when 6941 => read_data_o <= x"0000";
when 6942 => read_data_o <= x"0000";
when 6943 => read_data_o <= x"0000";
when 6944 => read_data_o <= x"0000";
when 6945 => read_data_o <= x"0000";
when 6946 => read_data_o <= x"0000";
when 6947 => read_data_o <= x"0000";
when 6948 => read_data_o <= x"0000";
when 6949 => read_data_o <= x"0000";
when 6950 => read_data_o <= x"0000";
when 6951 => read_data_o <= x"0000";
when 6952 => read_data_o <= x"0000";
when 6953 => read_data_o <= x"0000";
when 6954 => read_data_o <= x"0000";
when 6955 => read_data_o <= x"0000";
when 6956 => read_data_o <= x"0000";
when 6957 => read_data_o <= x"0000";
when 6958 => read_data_o <= x"0000";
when 6959 => read_data_o <= x"0000";
when 6960 => read_data_o <= x"0000";
when 6961 => read_data_o <= x"0000";
when 6962 => read_data_o <= x"0000";
when 6963 => read_data_o <= x"0000";
when 6964 => read_data_o <= x"0000";
when 6965 => read_data_o <= x"0000";
when 6966 => read_data_o <= x"0000";
when 6967 => read_data_o <= x"0000";
when 6968 => read_data_o <= x"0000";
when 6969 => read_data_o <= x"0000";
when 6970 => read_data_o <= x"0000";
when 6971 => read_data_o <= x"0000";
when 6972 => read_data_o <= x"0000";
when 6973 => read_data_o <= x"0000";
when 6974 => read_data_o <= x"0000";
when 6975 => read_data_o <= x"0000";
when 6976 => read_data_o <= x"0000";
when 6977 => read_data_o <= x"0000";
when 6978 => read_data_o <= x"0000";
when 6979 => read_data_o <= x"0000";
when 6980 => read_data_o <= x"0000";
when 6981 => read_data_o <= x"0000";
when 6982 => read_data_o <= x"0000";
when 6983 => read_data_o <= x"0000";
when 6984 => read_data_o <= x"0000";
when 6985 => read_data_o <= x"0000";
when 6986 => read_data_o <= x"0000";
when 6987 => read_data_o <= x"0000";
when 6988 => read_data_o <= x"0000";
when 6989 => read_data_o <= x"0000";
when 6990 => read_data_o <= x"0000";
when 6991 => read_data_o <= x"0000";
when 6992 => read_data_o <= x"0000";
when 6993 => read_data_o <= x"0000";
when 6994 => read_data_o <= x"0000";
when 6995 => read_data_o <= x"0000";
when 6996 => read_data_o <= x"0000";
when 6997 => read_data_o <= x"0000";
when 6998 => read_data_o <= x"0000";
when 6999 => read_data_o <= x"0000";
when 7000 => read_data_o <= x"0000";
when 7001 => read_data_o <= x"0000";
when 7002 => read_data_o <= x"0000";
when 7003 => read_data_o <= x"0000";
when 7004 => read_data_o <= x"0000";
when 7005 => read_data_o <= x"0000";
when 7006 => read_data_o <= x"0000";
when 7007 => read_data_o <= x"0000";
when 7008 => read_data_o <= x"0000";
when 7009 => read_data_o <= x"0000";
when 7010 => read_data_o <= x"0000";
when 7011 => read_data_o <= x"0000";
when 7012 => read_data_o <= x"d770";
when 7013 => read_data_o <= x"041a";
when 7014 => read_data_o <= x"0000";
when 7015 => read_data_o <= x"0000";
when 7016 => read_data_o <= x"001d";
when 7017 => read_data_o <= x"0000";
when 7018 => read_data_o <= x"0000";
when 7019 => read_data_o <= x"0000";
when 7020 => read_data_o <= x"0000";
when 7021 => read_data_o <= x"0000";
when 7022 => read_data_o <= x"0000";
when 7023 => read_data_o <= x"0000";
when 7024 => read_data_o <= x"0000";
when 7025 => read_data_o <= x"0000";
when 7026 => read_data_o <= x"0000";
when 7027 => read_data_o <= x"0000";
when 7028 => read_data_o <= x"0000";
when 7029 => read_data_o <= x"0000";
when 7030 => read_data_o <= x"0000";
when 7031 => read_data_o <= x"0000";
when 7032 => read_data_o <= x"0000";
when 7033 => read_data_o <= x"0000";
when 7034 => read_data_o <= x"0000";
when 7035 => read_data_o <= x"0000";
when 7036 => read_data_o <= x"0000";
when 7037 => read_data_o <= x"0000";
when 7038 => read_data_o <= x"0000";
when 7039 => read_data_o <= x"0000";
when 7040 => read_data_o <= x"0000";
when 7041 => read_data_o <= x"0000";
when 7042 => read_data_o <= x"0000";
when 7043 => read_data_o <= x"0000";
when 7044 => read_data_o <= x"0000";
when 7045 => read_data_o <= x"0000";
when 7046 => read_data_o <= x"0000";
when 7047 => read_data_o <= x"0000";
when 7048 => read_data_o <= x"0000";
when 7049 => read_data_o <= x"0000";
when 7050 => read_data_o <= x"0000";
when 7051 => read_data_o <= x"0000";
when 7052 => read_data_o <= x"0000";
when 7053 => read_data_o <= x"0000";
when 7054 => read_data_o <= x"0000";
when 7055 => read_data_o <= x"0000";
when 7056 => read_data_o <= x"0000";
when 7057 => read_data_o <= x"0000";
when 7058 => read_data_o <= x"0000";
when 7059 => read_data_o <= x"0000";
when 7060 => read_data_o <= x"0000";
when 7061 => read_data_o <= x"0000";
when 7062 => read_data_o <= x"0000";
when 7063 => read_data_o <= x"0000";
when 7064 => read_data_o <= x"0000";
when 7065 => read_data_o <= x"0000";
when 7066 => read_data_o <= x"0000";
when 7067 => read_data_o <= x"0000";
when 7068 => read_data_o <= x"0000";
when 7069 => read_data_o <= x"0000";
when 7070 => read_data_o <= x"0000";
when 7071 => read_data_o <= x"0000";
when 7072 => read_data_o <= x"0000";
when 7073 => read_data_o <= x"0000";
when 7074 => read_data_o <= x"0000";
when 7075 => read_data_o <= x"0000";
when 7076 => read_data_o <= x"0000";
when 7077 => read_data_o <= x"0000";
when 7078 => read_data_o <= x"0000";
when 7079 => read_data_o <= x"0000";
when 7080 => read_data_o <= x"0000";
when 7081 => read_data_o <= x"0000";
when 7082 => read_data_o <= x"0000";
when 7083 => read_data_o <= x"0000";
when 7084 => read_data_o <= x"0000";
when 7085 => read_data_o <= x"0000";
when 7086 => read_data_o <= x"0000";
when 7087 => read_data_o <= x"0000";
when 7088 => read_data_o <= x"0000";
when 7089 => read_data_o <= x"0000";
when 7090 => read_data_o <= x"0000";
when 7091 => read_data_o <= x"0000";
when 7092 => read_data_o <= x"d770";
when 7093 => read_data_o <= x"041a";
when 7094 => read_data_o <= x"0000";
when 7095 => read_data_o <= x"0000";
when 7096 => read_data_o <= x"001e";
when 7097 => read_data_o <= x"0000";
when 7098 => read_data_o <= x"0000";
when 7099 => read_data_o <= x"0000";
when 7100 => read_data_o <= x"0000";
when 7101 => read_data_o <= x"0000";
when 7102 => read_data_o <= x"d600";
when 7103 => read_data_o <= x"69be";
when 7104 => read_data_o <= x"0000";
when 7105 => read_data_o <= x"0000";
when 7106 => read_data_o <= x"0000";
when 7107 => read_data_o <= x"0000";
when 7108 => read_data_o <= x"0000";
when 7109 => read_data_o <= x"0000";
when 7110 => read_data_o <= x"0000";
when 7111 => read_data_o <= x"0000";
when 7112 => read_data_o <= x"0000";
when 7113 => read_data_o <= x"0000";
when 7114 => read_data_o <= x"0000";
when 7115 => read_data_o <= x"0000";
when 7116 => read_data_o <= x"0000";
when 7117 => read_data_o <= x"0000";
when 7118 => read_data_o <= x"0000";
when 7119 => read_data_o <= x"0000";
when 7120 => read_data_o <= x"0000";
when 7121 => read_data_o <= x"0000";
when 7122 => read_data_o <= x"0000";
when 7123 => read_data_o <= x"0000";
when 7124 => read_data_o <= x"0000";
when 7125 => read_data_o <= x"0000";
when 7126 => read_data_o <= x"0000";
when 7127 => read_data_o <= x"0000";
when 7128 => read_data_o <= x"0000";
when 7129 => read_data_o <= x"0000";
when 7130 => read_data_o <= x"0000";
when 7131 => read_data_o <= x"0000";
when 7132 => read_data_o <= x"0000";
when 7133 => read_data_o <= x"0000";
when 7134 => read_data_o <= x"0000";
when 7135 => read_data_o <= x"0000";
when 7136 => read_data_o <= x"0000";
when 7137 => read_data_o <= x"0000";
when 7138 => read_data_o <= x"0000";
when 7139 => read_data_o <= x"0000";
when 7140 => read_data_o <= x"0000";
when 7141 => read_data_o <= x"0000";
when 7142 => read_data_o <= x"0000";
when 7143 => read_data_o <= x"0000";
when 7144 => read_data_o <= x"0000";
when 7145 => read_data_o <= x"0000";
when 7146 => read_data_o <= x"0000";
when 7147 => read_data_o <= x"0000";
when 7148 => read_data_o <= x"0000";
when 7149 => read_data_o <= x"0000";
when 7150 => read_data_o <= x"0000";
when 7151 => read_data_o <= x"0000";
when 7152 => read_data_o <= x"0000";
when 7153 => read_data_o <= x"0000";
when 7154 => read_data_o <= x"0000";
when 7155 => read_data_o <= x"0000";
when 7156 => read_data_o <= x"0000";
when 7157 => read_data_o <= x"0000";
when 7158 => read_data_o <= x"0000";
when 7159 => read_data_o <= x"0000";
when 7160 => read_data_o <= x"0000";
when 7161 => read_data_o <= x"0000";
when 7162 => read_data_o <= x"0000";
when 7163 => read_data_o <= x"0000";
when 7164 => read_data_o <= x"0000";
when 7165 => read_data_o <= x"0000";
when 7166 => read_data_o <= x"0000";
when 7167 => read_data_o <= x"0000";
when 7168 => read_data_o <= x"0000";
when 7169 => read_data_o <= x"0000";
when 7170 => read_data_o <= x"5f63";
when 7171 => read_data_o <= x"7375";
when 7172 => read_data_o <= x"d770";
when 7173 => read_data_o <= x"041a";
when 7174 => read_data_o <= x"0000";
when 7175 => read_data_o <= x"0000";
when 7176 => read_data_o <= x"001f";
when 7177 => read_data_o <= x"0000";
when 7178 => read_data_o <= x"0000";
when 7179 => read_data_o <= x"0000";
when 7180 => read_data_o <= x"0000";
when 7181 => read_data_o <= x"0000";
when 7182 => read_data_o <= x"0000";
when 7183 => read_data_o <= x"0000";
when 7184 => read_data_o <= x"0000";
when 7185 => read_data_o <= x"0000";
when 7186 => read_data_o <= x"0000";
when 7187 => read_data_o <= x"0000";
when 7188 => read_data_o <= x"0000";
when 7189 => read_data_o <= x"0000";
when 7190 => read_data_o <= x"0000";
when 7191 => read_data_o <= x"0000";
when 7192 => read_data_o <= x"0000";
when 7193 => read_data_o <= x"0000";
when 7194 => read_data_o <= x"0000";
when 7195 => read_data_o <= x"0000";
when 7196 => read_data_o <= x"0000";
when 7197 => read_data_o <= x"0000";
when 7198 => read_data_o <= x"0000";
when 7199 => read_data_o <= x"0000";
when 7200 => read_data_o <= x"0000";
when 7201 => read_data_o <= x"0000";
when 7202 => read_data_o <= x"0000";
when 7203 => read_data_o <= x"0000";
when 7204 => read_data_o <= x"0000";
when 7205 => read_data_o <= x"0000";
when 7206 => read_data_o <= x"0000";
when 7207 => read_data_o <= x"0000";
when 7208 => read_data_o <= x"0000";
when 7209 => read_data_o <= x"0000";
when 7210 => read_data_o <= x"0000";
when 7211 => read_data_o <= x"0000";
when 7212 => read_data_o <= x"0000";
when 7213 => read_data_o <= x"0000";
when 7214 => read_data_o <= x"0000";
when 7215 => read_data_o <= x"0000";
when 7216 => read_data_o <= x"0000";
when 7217 => read_data_o <= x"0000";
when 7218 => read_data_o <= x"0000";
when 7219 => read_data_o <= x"0000";
when 7220 => read_data_o <= x"0000";
when 7221 => read_data_o <= x"0000";
when 7222 => read_data_o <= x"0000";
when 7223 => read_data_o <= x"0000";
when 7224 => read_data_o <= x"0000";
when 7225 => read_data_o <= x"0000";
when 7226 => read_data_o <= x"0000";
when 7227 => read_data_o <= x"0000";
when 7228 => read_data_o <= x"0000";
when 7229 => read_data_o <= x"0000";
when 7230 => read_data_o <= x"0000";
when 7231 => read_data_o <= x"0000";
when 7232 => read_data_o <= x"0000";
when 7233 => read_data_o <= x"0000";
when 7234 => read_data_o <= x"0000";
when 7235 => read_data_o <= x"0000";
when 7236 => read_data_o <= x"0000";
when 7237 => read_data_o <= x"0000";
when 7238 => read_data_o <= x"0000";
when 7239 => read_data_o <= x"0000";
when 7240 => read_data_o <= x"0000";
when 7241 => read_data_o <= x"0000";
when 7242 => read_data_o <= x"0000";
when 7243 => read_data_o <= x"0000";
when 7244 => read_data_o <= x"0000";
when 7245 => read_data_o <= x"0000";
when 7246 => read_data_o <= x"0000";
when 7247 => read_data_o <= x"0000";
when 7248 => read_data_o <= x"0000";
when 7249 => read_data_o <= x"0000";
when 7250 => read_data_o <= x"0000";
when 7251 => read_data_o <= x"0000";
when 7252 => read_data_o <= x"d770";
when 7253 => read_data_o <= x"041a";
when 7254 => read_data_o <= x"0000";
when 7255 => read_data_o <= x"0000";
when 7256 => read_data_o <= x"0020";
when 7257 => read_data_o <= x"0000";
when 7258 => read_data_o <= x"0000";
when 7259 => read_data_o <= x"0000";
when 7260 => read_data_o <= x"0000";
when 7261 => read_data_o <= x"0000";
when 7262 => read_data_o <= x"0000";
when 7263 => read_data_o <= x"0000";
when 7264 => read_data_o <= x"0000";
when 7265 => read_data_o <= x"0000";
when 7266 => read_data_o <= x"0000";
when 7267 => read_data_o <= x"0000";
when 7268 => read_data_o <= x"0000";
when 7269 => read_data_o <= x"0000";
when 7270 => read_data_o <= x"0000";
when 7271 => read_data_o <= x"0000";
when 7272 => read_data_o <= x"0000";
when 7273 => read_data_o <= x"0000";
when 7274 => read_data_o <= x"0000";
when 7275 => read_data_o <= x"0000";
when 7276 => read_data_o <= x"0000";
when 7277 => read_data_o <= x"0000";
when 7278 => read_data_o <= x"0000";
when 7279 => read_data_o <= x"0000";
when 7280 => read_data_o <= x"0000";
when 7281 => read_data_o <= x"0000";
when 7282 => read_data_o <= x"0000";
when 7283 => read_data_o <= x"0000";
when 7284 => read_data_o <= x"0000";
when 7285 => read_data_o <= x"0000";
when 7286 => read_data_o <= x"0000";
when 7287 => read_data_o <= x"0000";
when 7288 => read_data_o <= x"0000";
when 7289 => read_data_o <= x"0000";
when 7290 => read_data_o <= x"0000";
when 7291 => read_data_o <= x"0000";
when 7292 => read_data_o <= x"0000";
when 7293 => read_data_o <= x"0000";
when 7294 => read_data_o <= x"0000";
when 7295 => read_data_o <= x"0000";
when 7296 => read_data_o <= x"0000";
when 7297 => read_data_o <= x"0000";
when 7298 => read_data_o <= x"0000";
when 7299 => read_data_o <= x"0000";
when 7300 => read_data_o <= x"0000";
when 7301 => read_data_o <= x"0000";
when 7302 => read_data_o <= x"0000";
when 7303 => read_data_o <= x"0000";
when 7304 => read_data_o <= x"0000";
when 7305 => read_data_o <= x"0000";
when 7306 => read_data_o <= x"0000";
when 7307 => read_data_o <= x"0000";
when 7308 => read_data_o <= x"0000";
when 7309 => read_data_o <= x"0000";
when 7310 => read_data_o <= x"0000";
when 7311 => read_data_o <= x"0000";
when 7312 => read_data_o <= x"0000";
when 7313 => read_data_o <= x"0000";
when 7314 => read_data_o <= x"0000";
when 7315 => read_data_o <= x"0000";
when 7316 => read_data_o <= x"0000";
when 7317 => read_data_o <= x"0000";
when 7318 => read_data_o <= x"0000";
when 7319 => read_data_o <= x"0000";
when 7320 => read_data_o <= x"0000";
when 7321 => read_data_o <= x"0000";
when 7322 => read_data_o <= x"0000";
when 7323 => read_data_o <= x"0000";
when 7324 => read_data_o <= x"0000";
when 7325 => read_data_o <= x"0000";
when 7326 => read_data_o <= x"0000";
when 7327 => read_data_o <= x"0000";
when 7328 => read_data_o <= x"0000";
when 7329 => read_data_o <= x"0000";
when 7330 => read_data_o <= x"0000";
when 7331 => read_data_o <= x"0000";
when 7332 => read_data_o <= x"d770";
when 7333 => read_data_o <= x"041a";
when 7334 => read_data_o <= x"0000";
when 7335 => read_data_o <= x"0000";
when 7336 => read_data_o <= x"0021";
when 7337 => read_data_o <= x"0000";
when 7338 => read_data_o <= x"0000";
when 7339 => read_data_o <= x"0000";
when 7340 => read_data_o <= x"0000";
when 7341 => read_data_o <= x"0000";
when 7342 => read_data_o <= x"ff00";
when 7343 => read_data_o <= x"ffff";
when 7344 => read_data_o <= x"0000";
when 7345 => read_data_o <= x"0000";
when 7346 => read_data_o <= x"0000";
when 7347 => read_data_o <= x"0000";
when 7348 => read_data_o <= x"0000";
when 7349 => read_data_o <= x"0000";
when 7350 => read_data_o <= x"0000";
when 7351 => read_data_o <= x"0000";
when 7352 => read_data_o <= x"0000";
when 7353 => read_data_o <= x"0000";
when 7354 => read_data_o <= x"0000";
when 7355 => read_data_o <= x"0000";
when 7356 => read_data_o <= x"0000";
when 7357 => read_data_o <= x"0000";
when 7358 => read_data_o <= x"0000";
when 7359 => read_data_o <= x"0000";
when 7360 => read_data_o <= x"0000";
when 7361 => read_data_o <= x"0000";
when 7362 => read_data_o <= x"0000";
when 7363 => read_data_o <= x"0000";
when 7364 => read_data_o <= x"0000";
when 7365 => read_data_o <= x"0000";
when 7366 => read_data_o <= x"0000";
when 7367 => read_data_o <= x"0000";
when 7368 => read_data_o <= x"0000";
when 7369 => read_data_o <= x"0000";
when 7370 => read_data_o <= x"0000";
when 7371 => read_data_o <= x"0000";
when 7372 => read_data_o <= x"0000";
when 7373 => read_data_o <= x"0000";
when 7374 => read_data_o <= x"0000";
when 7375 => read_data_o <= x"0000";
when 7376 => read_data_o <= x"0000";
when 7377 => read_data_o <= x"0000";
when 7378 => read_data_o <= x"0000";
when 7379 => read_data_o <= x"0000";
when 7380 => read_data_o <= x"0000";
when 7381 => read_data_o <= x"0000";
when 7382 => read_data_o <= x"0000";
when 7383 => read_data_o <= x"0000";
when 7384 => read_data_o <= x"0000";
when 7385 => read_data_o <= x"0000";
when 7386 => read_data_o <= x"0000";
when 7387 => read_data_o <= x"0000";
when 7388 => read_data_o <= x"0000";
when 7389 => read_data_o <= x"0000";
when 7390 => read_data_o <= x"0000";
when 7391 => read_data_o <= x"0000";
when 7392 => read_data_o <= x"0000";
when 7393 => read_data_o <= x"0000";
when 7394 => read_data_o <= x"0000";
when 7395 => read_data_o <= x"0000";
when 7396 => read_data_o <= x"0000";
when 7397 => read_data_o <= x"0000";
when 7398 => read_data_o <= x"0000";
when 7399 => read_data_o <= x"0000";
when 7400 => read_data_o <= x"0000";
when 7401 => read_data_o <= x"0000";
when 7402 => read_data_o <= x"0000";
when 7403 => read_data_o <= x"0000";
when 7404 => read_data_o <= x"0000";
when 7405 => read_data_o <= x"0000";
when 7406 => read_data_o <= x"0000";
when 7407 => read_data_o <= x"0000";
when 7408 => read_data_o <= x"0000";
when 7409 => read_data_o <= x"0000";
when 7410 => read_data_o <= x"0000";
when 7411 => read_data_o <= x"0000";
when 7412 => read_data_o <= x"d770";
when 7413 => read_data_o <= x"041a";
when 7414 => read_data_o <= x"0000";
when 7415 => read_data_o <= x"0000";
when 7416 => read_data_o <= x"0022";
when 7417 => read_data_o <= x"0000";
when 7418 => read_data_o <= x"0000";
when 7419 => read_data_o <= x"0000";
when 7420 => read_data_o <= x"0000";
when 7421 => read_data_o <= x"0000";
when 7422 => read_data_o <= x"4700";
when 7423 => read_data_o <= x"976e";
when 7424 => read_data_o <= x"0000";
when 7425 => read_data_o <= x"0000";
when 7426 => read_data_o <= x"0000";
when 7427 => read_data_o <= x"0000";
when 7428 => read_data_o <= x"0000";
when 7429 => read_data_o <= x"0000";
when 7430 => read_data_o <= x"0000";
when 7431 => read_data_o <= x"0000";
when 7432 => read_data_o <= x"0000";
when 7433 => read_data_o <= x"0000";
when 7434 => read_data_o <= x"0000";
when 7435 => read_data_o <= x"0000";
when 7436 => read_data_o <= x"0000";
when 7437 => read_data_o <= x"0000";
when 7438 => read_data_o <= x"0000";
when 7439 => read_data_o <= x"0000";
when 7440 => read_data_o <= x"0000";
when 7441 => read_data_o <= x"0000";
when 7442 => read_data_o <= x"0000";
when 7443 => read_data_o <= x"0000";
when 7444 => read_data_o <= x"0000";
when 7445 => read_data_o <= x"0000";
when 7446 => read_data_o <= x"0000";
when 7447 => read_data_o <= x"0000";
when 7448 => read_data_o <= x"0000";
when 7449 => read_data_o <= x"0000";
when 7450 => read_data_o <= x"0000";
when 7451 => read_data_o <= x"0000";
when 7452 => read_data_o <= x"0000";
when 7453 => read_data_o <= x"0000";
when 7454 => read_data_o <= x"0000";
when 7455 => read_data_o <= x"0000";
when 7456 => read_data_o <= x"0000";
when 7457 => read_data_o <= x"0000";
when 7458 => read_data_o <= x"0000";
when 7459 => read_data_o <= x"0000";
when 7460 => read_data_o <= x"0000";
when 7461 => read_data_o <= x"0000";
when 7462 => read_data_o <= x"0000";
when 7463 => read_data_o <= x"0000";
when 7464 => read_data_o <= x"0000";
when 7465 => read_data_o <= x"0000";
when 7466 => read_data_o <= x"0000";
when 7467 => read_data_o <= x"0000";
when 7468 => read_data_o <= x"0000";
when 7469 => read_data_o <= x"0000";
when 7470 => read_data_o <= x"0000";
when 7471 => read_data_o <= x"0000";
when 7472 => read_data_o <= x"0000";
when 7473 => read_data_o <= x"0000";
when 7474 => read_data_o <= x"0000";
when 7475 => read_data_o <= x"0000";
when 7476 => read_data_o <= x"0000";
when 7477 => read_data_o <= x"0000";
when 7478 => read_data_o <= x"0000";
when 7479 => read_data_o <= x"0000";
when 7480 => read_data_o <= x"0000";
when 7481 => read_data_o <= x"0000";
when 7482 => read_data_o <= x"0000";
when 7483 => read_data_o <= x"0000";
when 7484 => read_data_o <= x"0000";
when 7485 => read_data_o <= x"0000";
when 7486 => read_data_o <= x"0000";
when 7487 => read_data_o <= x"0000";
when 7488 => read_data_o <= x"0000";
when 7489 => read_data_o <= x"0000";
when 7490 => read_data_o <= x"0000";
when 7491 => read_data_o <= x"0000";
when 7492 => read_data_o <= x"d770";
when 7493 => read_data_o <= x"041a";
when 7494 => read_data_o <= x"0000";
when 7495 => read_data_o <= x"0000";
when 7496 => read_data_o <= x"0023";
when 7497 => read_data_o <= x"0000";
when 7498 => read_data_o <= x"0000";
when 7499 => read_data_o <= x"0000";
when 7500 => read_data_o <= x"0000";
when 7501 => read_data_o <= x"0000";
when 7502 => read_data_o <= x"0000";
when 7503 => read_data_o <= x"0000";
when 7504 => read_data_o <= x"0000";
when 7505 => read_data_o <= x"0000";
when 7506 => read_data_o <= x"0000";
when 7507 => read_data_o <= x"0000";
when 7508 => read_data_o <= x"0000";
when 7509 => read_data_o <= x"0000";
when 7510 => read_data_o <= x"0000";
when 7511 => read_data_o <= x"0000";
when 7512 => read_data_o <= x"0000";
when 7513 => read_data_o <= x"0000";
when 7514 => read_data_o <= x"0000";
when 7515 => read_data_o <= x"0000";
when 7516 => read_data_o <= x"0000";
when 7517 => read_data_o <= x"0000";
when 7518 => read_data_o <= x"0000";
when 7519 => read_data_o <= x"0000";
when 7520 => read_data_o <= x"0000";
when 7521 => read_data_o <= x"0000";
when 7522 => read_data_o <= x"0000";
when 7523 => read_data_o <= x"0000";
when 7524 => read_data_o <= x"0000";
when 7525 => read_data_o <= x"0000";
when 7526 => read_data_o <= x"0000";
when 7527 => read_data_o <= x"0000";
when 7528 => read_data_o <= x"0000";
when 7529 => read_data_o <= x"0000";
when 7530 => read_data_o <= x"0000";
when 7531 => read_data_o <= x"0000";
when 7532 => read_data_o <= x"0000";
when 7533 => read_data_o <= x"0000";
when 7534 => read_data_o <= x"0000";
when 7535 => read_data_o <= x"0000";
when 7536 => read_data_o <= x"0000";
when 7537 => read_data_o <= x"0000";
when 7538 => read_data_o <= x"0000";
when 7539 => read_data_o <= x"0000";
when 7540 => read_data_o <= x"0000";
when 7541 => read_data_o <= x"0000";
when 7542 => read_data_o <= x"0000";
when 7543 => read_data_o <= x"0000";
when 7544 => read_data_o <= x"0000";
when 7545 => read_data_o <= x"0000";
when 7546 => read_data_o <= x"0000";
when 7547 => read_data_o <= x"0000";
when 7548 => read_data_o <= x"0000";
when 7549 => read_data_o <= x"0000";
when 7550 => read_data_o <= x"0000";
when 7551 => read_data_o <= x"0000";
when 7552 => read_data_o <= x"0000";
when 7553 => read_data_o <= x"0000";
when 7554 => read_data_o <= x"0000";
when 7555 => read_data_o <= x"0000";
when 7556 => read_data_o <= x"0000";
when 7557 => read_data_o <= x"0000";
when 7558 => read_data_o <= x"0000";
when 7559 => read_data_o <= x"0000";
when 7560 => read_data_o <= x"0000";
when 7561 => read_data_o <= x"0000";
when 7562 => read_data_o <= x"0000";
when 7563 => read_data_o <= x"0000";
when 7564 => read_data_o <= x"0000";
when 7565 => read_data_o <= x"0000";
when 7566 => read_data_o <= x"0000";
when 7567 => read_data_o <= x"0000";
when 7568 => read_data_o <= x"0000";
when 7569 => read_data_o <= x"0000";
when 7570 => read_data_o <= x"0000";
when 7571 => read_data_o <= x"0000";
when 7572 => read_data_o <= x"d770";
when 7573 => read_data_o <= x"041a";
when 7574 => read_data_o <= x"0000";
when 7575 => read_data_o <= x"0000";
when 7576 => read_data_o <= x"0024";
when 7577 => read_data_o <= x"0000";
when 7578 => read_data_o <= x"0000";
when 7579 => read_data_o <= x"0000";
when 7580 => read_data_o <= x"0000";
when 7581 => read_data_o <= x"0000";
when 7582 => read_data_o <= x"7f00";
when 7583 => read_data_o <= x"0000";
when 7584 => read_data_o <= x"0000";
when 7585 => read_data_o <= x"0000";
when 7586 => read_data_o <= x"0000";
when 7587 => read_data_o <= x"0000";
when 7588 => read_data_o <= x"0000";
when 7589 => read_data_o <= x"0000";
when 7590 => read_data_o <= x"0000";
when 7591 => read_data_o <= x"0000";
when 7592 => read_data_o <= x"0000";
when 7593 => read_data_o <= x"0000";
when 7594 => read_data_o <= x"0000";
when 7595 => read_data_o <= x"0000";
when 7596 => read_data_o <= x"0000";
when 7597 => read_data_o <= x"0000";
when 7598 => read_data_o <= x"0000";
when 7599 => read_data_o <= x"0000";
when 7600 => read_data_o <= x"0000";
when 7601 => read_data_o <= x"0000";
when 7602 => read_data_o <= x"0000";
when 7603 => read_data_o <= x"0000";
when 7604 => read_data_o <= x"0000";
when 7605 => read_data_o <= x"0000";
when 7606 => read_data_o <= x"0000";
when 7607 => read_data_o <= x"0000";
when 7608 => read_data_o <= x"0000";
when 7609 => read_data_o <= x"0000";
when 7610 => read_data_o <= x"0000";
when 7611 => read_data_o <= x"0000";
when 7612 => read_data_o <= x"0000";
when 7613 => read_data_o <= x"0000";
when 7614 => read_data_o <= x"0000";
when 7615 => read_data_o <= x"0000";
when 7616 => read_data_o <= x"0000";
when 7617 => read_data_o <= x"0000";
when 7618 => read_data_o <= x"0000";
when 7619 => read_data_o <= x"0000";
when 7620 => read_data_o <= x"0000";
when 7621 => read_data_o <= x"0000";
when 7622 => read_data_o <= x"0000";
when 7623 => read_data_o <= x"0000";
when 7624 => read_data_o <= x"0000";
when 7625 => read_data_o <= x"0000";
when 7626 => read_data_o <= x"0000";
when 7627 => read_data_o <= x"0000";
when 7628 => read_data_o <= x"0000";
when 7629 => read_data_o <= x"0000";
when 7630 => read_data_o <= x"0000";
when 7631 => read_data_o <= x"0000";
when 7632 => read_data_o <= x"0000";
when 7633 => read_data_o <= x"0000";
when 7634 => read_data_o <= x"0000";
when 7635 => read_data_o <= x"0000";
when 7636 => read_data_o <= x"0000";
when 7637 => read_data_o <= x"0000";
when 7638 => read_data_o <= x"0000";
when 7639 => read_data_o <= x"0000";
when 7640 => read_data_o <= x"0000";
when 7641 => read_data_o <= x"0000";
when 7642 => read_data_o <= x"0000";
when 7643 => read_data_o <= x"0000";
when 7644 => read_data_o <= x"0000";
when 7645 => read_data_o <= x"0000";
when 7646 => read_data_o <= x"0000";
when 7647 => read_data_o <= x"0000";
when 7648 => read_data_o <= x"0000";
when 7649 => read_data_o <= x"0000";
when 7650 => read_data_o <= x"0000";
when 7651 => read_data_o <= x"0000";
when 7652 => read_data_o <= x"d770";
when 7653 => read_data_o <= x"041a";
when 7654 => read_data_o <= x"0000";
when 7655 => read_data_o <= x"0000";
when 7656 => read_data_o <= x"0025";
when 7657 => read_data_o <= x"0000";
when 7658 => read_data_o <= x"0000";
when 7659 => read_data_o <= x"0000";
when 7660 => read_data_o <= x"0000";
when 7661 => read_data_o <= x"0000";
when 7662 => read_data_o <= x"0000";
when 7663 => read_data_o <= x"0000";
when 7664 => read_data_o <= x"0000";
when 7665 => read_data_o <= x"0000";
when 7666 => read_data_o <= x"0000";
when 7667 => read_data_o <= x"0000";
when 7668 => read_data_o <= x"0000";
when 7669 => read_data_o <= x"0000";
when 7670 => read_data_o <= x"0000";
when 7671 => read_data_o <= x"0000";
when 7672 => read_data_o <= x"0000";
when 7673 => read_data_o <= x"0000";
when 7674 => read_data_o <= x"0000";
when 7675 => read_data_o <= x"0000";
when 7676 => read_data_o <= x"0000";
when 7677 => read_data_o <= x"0000";
when 7678 => read_data_o <= x"0000";
when 7679 => read_data_o <= x"0000";
when 7680 => read_data_o <= x"0000";
when 7681 => read_data_o <= x"0000";
when 7682 => read_data_o <= x"0000";
when 7683 => read_data_o <= x"0000";
when 7684 => read_data_o <= x"0000";
when 7685 => read_data_o <= x"0000";
when 7686 => read_data_o <= x"0000";
when 7687 => read_data_o <= x"0000";
when 7688 => read_data_o <= x"0000";
when 7689 => read_data_o <= x"0000";
when 7690 => read_data_o <= x"0000";
when 7691 => read_data_o <= x"0000";
when 7692 => read_data_o <= x"0000";
when 7693 => read_data_o <= x"0000";
when 7694 => read_data_o <= x"0000";
when 7695 => read_data_o <= x"0000";
when 7696 => read_data_o <= x"0000";
when 7697 => read_data_o <= x"0000";
when 7698 => read_data_o <= x"0000";
when 7699 => read_data_o <= x"0000";
when 7700 => read_data_o <= x"0000";
when 7701 => read_data_o <= x"0000";
when 7702 => read_data_o <= x"0000";
when 7703 => read_data_o <= x"0000";
when 7704 => read_data_o <= x"0000";
when 7705 => read_data_o <= x"0000";
when 7706 => read_data_o <= x"0000";
when 7707 => read_data_o <= x"0000";
when 7708 => read_data_o <= x"0000";
when 7709 => read_data_o <= x"0000";
when 7710 => read_data_o <= x"0000";
when 7711 => read_data_o <= x"0000";
when 7712 => read_data_o <= x"0000";
when 7713 => read_data_o <= x"0000";
when 7714 => read_data_o <= x"0000";
when 7715 => read_data_o <= x"0000";
when 7716 => read_data_o <= x"0000";
when 7717 => read_data_o <= x"0000";
when 7718 => read_data_o <= x"0000";
when 7719 => read_data_o <= x"0000";
when 7720 => read_data_o <= x"0000";
when 7721 => read_data_o <= x"0000";
when 7722 => read_data_o <= x"0000";
when 7723 => read_data_o <= x"0000";
when 7724 => read_data_o <= x"0000";
when 7725 => read_data_o <= x"0000";
when 7726 => read_data_o <= x"0000";
when 7727 => read_data_o <= x"0000";
when 7728 => read_data_o <= x"0000";
when 7729 => read_data_o <= x"0000";
when 7730 => read_data_o <= x"0000";
when 7731 => read_data_o <= x"0000";
when 7732 => read_data_o <= x"d770";
when 7733 => read_data_o <= x"041a";
when 7734 => read_data_o <= x"0000";
when 7735 => read_data_o <= x"0000";
when 7736 => read_data_o <= x"0026";
when 7737 => read_data_o <= x"0000";
when 7738 => read_data_o <= x"0000";
when 7739 => read_data_o <= x"0000";
when 7740 => read_data_o <= x"0000";
when 7741 => read_data_o <= x"0000";
when 7742 => read_data_o <= x"0000";
when 7743 => read_data_o <= x"0000";
when 7744 => read_data_o <= x"0000";
when 7745 => read_data_o <= x"0000";
when 7746 => read_data_o <= x"0000";
when 7747 => read_data_o <= x"0000";
when 7748 => read_data_o <= x"0000";
when 7749 => read_data_o <= x"0000";
when 7750 => read_data_o <= x"0000";
when 7751 => read_data_o <= x"0000";
when 7752 => read_data_o <= x"0000";
when 7753 => read_data_o <= x"0000";
when 7754 => read_data_o <= x"0000";
when 7755 => read_data_o <= x"0000";
when 7756 => read_data_o <= x"0000";
when 7757 => read_data_o <= x"0000";
when 7758 => read_data_o <= x"0000";
when 7759 => read_data_o <= x"0000";
when 7760 => read_data_o <= x"0000";
when 7761 => read_data_o <= x"0000";
when 7762 => read_data_o <= x"0000";
when 7763 => read_data_o <= x"0000";
when 7764 => read_data_o <= x"0000";
when 7765 => read_data_o <= x"0000";
when 7766 => read_data_o <= x"0000";
when 7767 => read_data_o <= x"0000";
when 7768 => read_data_o <= x"0000";
when 7769 => read_data_o <= x"0000";
when 7770 => read_data_o <= x"0000";
when 7771 => read_data_o <= x"0000";
when 7772 => read_data_o <= x"0000";
when 7773 => read_data_o <= x"0000";
when 7774 => read_data_o <= x"0000";
when 7775 => read_data_o <= x"0000";
when 7776 => read_data_o <= x"0000";
when 7777 => read_data_o <= x"0000";
when 7778 => read_data_o <= x"0000";
when 7779 => read_data_o <= x"0000";
when 7780 => read_data_o <= x"0000";
when 7781 => read_data_o <= x"0000";
when 7782 => read_data_o <= x"0000";
when 7783 => read_data_o <= x"0000";
when 7784 => read_data_o <= x"0000";
when 7785 => read_data_o <= x"0000";
when 7786 => read_data_o <= x"0000";
when 7787 => read_data_o <= x"0000";
when 7788 => read_data_o <= x"0000";
when 7789 => read_data_o <= x"0000";
when 7790 => read_data_o <= x"0000";
when 7791 => read_data_o <= x"0000";
when 7792 => read_data_o <= x"0000";
when 7793 => read_data_o <= x"0000";
when 7794 => read_data_o <= x"0000";
when 7795 => read_data_o <= x"0000";
when 7796 => read_data_o <= x"0000";
when 7797 => read_data_o <= x"0000";
when 7798 => read_data_o <= x"0000";
when 7799 => read_data_o <= x"0000";
when 7800 => read_data_o <= x"0000";
when 7801 => read_data_o <= x"0000";
when 7802 => read_data_o <= x"0000";
when 7803 => read_data_o <= x"0000";
when 7804 => read_data_o <= x"0000";
when 7805 => read_data_o <= x"0000";
when 7806 => read_data_o <= x"0000";
when 7807 => read_data_o <= x"0000";
when 7808 => read_data_o <= x"0000";
when 7809 => read_data_o <= x"0000";
when 7810 => read_data_o <= x"0000";
when 7811 => read_data_o <= x"0000";
when 7812 => read_data_o <= x"d770";
when 7813 => read_data_o <= x"041a";
when 7814 => read_data_o <= x"0000";
when 7815 => read_data_o <= x"0000";
when 7816 => read_data_o <= x"0027";
when 7817 => read_data_o <= x"0000";
when 7818 => read_data_o <= x"0000";
when 7819 => read_data_o <= x"0000";
when 7820 => read_data_o <= x"0000";
when 7821 => read_data_o <= x"0000";
when 7822 => read_data_o <= x"0000";
when 7823 => read_data_o <= x"0000";
when 7824 => read_data_o <= x"0000";
when 7825 => read_data_o <= x"0000";
when 7826 => read_data_o <= x"0000";
when 7827 => read_data_o <= x"0000";
when 7828 => read_data_o <= x"0000";
when 7829 => read_data_o <= x"0000";
when 7830 => read_data_o <= x"0000";
when 7831 => read_data_o <= x"0000";
when 7832 => read_data_o <= x"0000";
when 7833 => read_data_o <= x"0000";
when 7834 => read_data_o <= x"0000";
when 7835 => read_data_o <= x"0000";
when 7836 => read_data_o <= x"0000";
when 7837 => read_data_o <= x"0000";
when 7838 => read_data_o <= x"0000";
when 7839 => read_data_o <= x"0000";
when 7840 => read_data_o <= x"0000";
when 7841 => read_data_o <= x"0000";
when 7842 => read_data_o <= x"0000";
when 7843 => read_data_o <= x"0000";
when 7844 => read_data_o <= x"0000";
when 7845 => read_data_o <= x"0000";
when 7846 => read_data_o <= x"0000";
when 7847 => read_data_o <= x"0000";
when 7848 => read_data_o <= x"0000";
when 7849 => read_data_o <= x"0000";
when 7850 => read_data_o <= x"0000";
when 7851 => read_data_o <= x"0000";
when 7852 => read_data_o <= x"0000";
when 7853 => read_data_o <= x"0000";
when 7854 => read_data_o <= x"0000";
when 7855 => read_data_o <= x"0000";
when 7856 => read_data_o <= x"0000";
when 7857 => read_data_o <= x"0000";
when 7858 => read_data_o <= x"0000";
when 7859 => read_data_o <= x"0000";
when 7860 => read_data_o <= x"0000";
when 7861 => read_data_o <= x"0000";
when 7862 => read_data_o <= x"0000";
when 7863 => read_data_o <= x"0000";
when 7864 => read_data_o <= x"0000";
when 7865 => read_data_o <= x"0000";
when 7866 => read_data_o <= x"0000";
when 7867 => read_data_o <= x"0000";
when 7868 => read_data_o <= x"0000";
when 7869 => read_data_o <= x"0000";
when 7870 => read_data_o <= x"0000";
when 7871 => read_data_o <= x"0000";
when 7872 => read_data_o <= x"0000";
when 7873 => read_data_o <= x"0000";
when 7874 => read_data_o <= x"0000";
when 7875 => read_data_o <= x"0000";
when 7876 => read_data_o <= x"0000";
when 7877 => read_data_o <= x"0000";
when 7878 => read_data_o <= x"0000";
when 7879 => read_data_o <= x"0000";
when 7880 => read_data_o <= x"0000";
when 7881 => read_data_o <= x"0000";
when 7882 => read_data_o <= x"0000";
when 7883 => read_data_o <= x"0000";
when 7884 => read_data_o <= x"0000";
when 7885 => read_data_o <= x"0000";
when 7886 => read_data_o <= x"0000";
when 7887 => read_data_o <= x"0000";
when 7888 => read_data_o <= x"0000";
when 7889 => read_data_o <= x"0000";
when 7890 => read_data_o <= x"6f72";
when 7891 => read_data_o <= x"006c";
when 7892 => read_data_o <= x"d770";
when 7893 => read_data_o <= x"041a";
when 7894 => read_data_o <= x"0000";
when 7895 => read_data_o <= x"0000";
when 7896 => read_data_o <= x"0028";
when 7897 => read_data_o <= x"0000";
when 7898 => read_data_o <= x"0000";
when 7899 => read_data_o <= x"0000";
when 7900 => read_data_o <= x"0000";
when 7901 => read_data_o <= x"0000";
when 7902 => read_data_o <= x"0000";
when 7903 => read_data_o <= x"0000";
when 7904 => read_data_o <= x"0000";
when 7905 => read_data_o <= x"0000";
when 7906 => read_data_o <= x"0000";
when 7907 => read_data_o <= x"0000";
when 7908 => read_data_o <= x"0000";
when 7909 => read_data_o <= x"0000";
when 7910 => read_data_o <= x"0000";
when 7911 => read_data_o <= x"0000";
when 7912 => read_data_o <= x"0000";
when 7913 => read_data_o <= x"0000";
when 7914 => read_data_o <= x"0000";
when 7915 => read_data_o <= x"0000";
when 7916 => read_data_o <= x"0000";
when 7917 => read_data_o <= x"0000";
when 7918 => read_data_o <= x"0000";
when 7919 => read_data_o <= x"0000";
when 7920 => read_data_o <= x"0000";
when 7921 => read_data_o <= x"0000";
when 7922 => read_data_o <= x"0000";
when 7923 => read_data_o <= x"0000";
when 7924 => read_data_o <= x"0000";
when 7925 => read_data_o <= x"0000";
when 7926 => read_data_o <= x"0000";
when 7927 => read_data_o <= x"0000";
when 7928 => read_data_o <= x"0000";
when 7929 => read_data_o <= x"0000";
when 7930 => read_data_o <= x"0000";
when 7931 => read_data_o <= x"0000";
when 7932 => read_data_o <= x"0000";
when 7933 => read_data_o <= x"0000";
when 7934 => read_data_o <= x"0000";
when 7935 => read_data_o <= x"0000";
when 7936 => read_data_o <= x"0000";
when 7937 => read_data_o <= x"0000";
when 7938 => read_data_o <= x"0000";
when 7939 => read_data_o <= x"0000";
when 7940 => read_data_o <= x"0000";
when 7941 => read_data_o <= x"0000";
when 7942 => read_data_o <= x"0000";
when 7943 => read_data_o <= x"0000";
when 7944 => read_data_o <= x"0000";
when 7945 => read_data_o <= x"0000";
when 7946 => read_data_o <= x"0000";
when 7947 => read_data_o <= x"0000";
when 7948 => read_data_o <= x"0000";
when 7949 => read_data_o <= x"0000";
when 7950 => read_data_o <= x"0000";
when 7951 => read_data_o <= x"0000";
when 7952 => read_data_o <= x"0000";
when 7953 => read_data_o <= x"0000";
when 7954 => read_data_o <= x"0000";
when 7955 => read_data_o <= x"0000";
when 7956 => read_data_o <= x"0000";
when 7957 => read_data_o <= x"0000";
when 7958 => read_data_o <= x"0000";
when 7959 => read_data_o <= x"0000";
when 7960 => read_data_o <= x"0000";
when 7961 => read_data_o <= x"0000";
when 7962 => read_data_o <= x"0000";
when 7963 => read_data_o <= x"0000";
when 7964 => read_data_o <= x"0000";
when 7965 => read_data_o <= x"0000";
when 7966 => read_data_o <= x"0000";
when 7967 => read_data_o <= x"0000";
when 7968 => read_data_o <= x"0000";
when 7969 => read_data_o <= x"0000";
when 7970 => read_data_o <= x"0000";
when 7971 => read_data_o <= x"0000";
when 7972 => read_data_o <= x"d770";
when 7973 => read_data_o <= x"041a";
when 7974 => read_data_o <= x"0000";
when 7975 => read_data_o <= x"0000";
when 7976 => read_data_o <= x"0029";
when 7977 => read_data_o <= x"0000";
when 7978 => read_data_o <= x"0000";
when 7979 => read_data_o <= x"0000";
when 7980 => read_data_o <= x"0000";
when 7981 => read_data_o <= x"0000";
when 7982 => read_data_o <= x"0000";
when 7983 => read_data_o <= x"0000";
when 7984 => read_data_o <= x"0000";
when 7985 => read_data_o <= x"0000";
when 7986 => read_data_o <= x"0000";
when 7987 => read_data_o <= x"0000";
when 7988 => read_data_o <= x"0000";
when 7989 => read_data_o <= x"0000";
when 7990 => read_data_o <= x"0000";
when 7991 => read_data_o <= x"0000";
when 7992 => read_data_o <= x"0000";
when 7993 => read_data_o <= x"0000";
when 7994 => read_data_o <= x"0000";
when 7995 => read_data_o <= x"0000";
when 7996 => read_data_o <= x"0000";
when 7997 => read_data_o <= x"0000";
when 7998 => read_data_o <= x"0000";
when 7999 => read_data_o <= x"0000";
when 8000 => read_data_o <= x"0000";
when 8001 => read_data_o <= x"0000";
when 8002 => read_data_o <= x"0000";
when 8003 => read_data_o <= x"0000";
when 8004 => read_data_o <= x"0000";
when 8005 => read_data_o <= x"0000";
when 8006 => read_data_o <= x"0000";
when 8007 => read_data_o <= x"0000";
when 8008 => read_data_o <= x"0000";
when 8009 => read_data_o <= x"0000";
when 8010 => read_data_o <= x"0000";
when 8011 => read_data_o <= x"0000";
when 8012 => read_data_o <= x"0000";
when 8013 => read_data_o <= x"0000";
when 8014 => read_data_o <= x"0000";
when 8015 => read_data_o <= x"0000";
when 8016 => read_data_o <= x"0000";
when 8017 => read_data_o <= x"0000";
when 8018 => read_data_o <= x"0000";
when 8019 => read_data_o <= x"0000";
when 8020 => read_data_o <= x"0000";
when 8021 => read_data_o <= x"0000";
when 8022 => read_data_o <= x"0000";
when 8023 => read_data_o <= x"0000";
when 8024 => read_data_o <= x"0000";
when 8025 => read_data_o <= x"0000";
when 8026 => read_data_o <= x"0000";
when 8027 => read_data_o <= x"0000";
when 8028 => read_data_o <= x"0000";
when 8029 => read_data_o <= x"0000";
when 8030 => read_data_o <= x"0000";
when 8031 => read_data_o <= x"0000";
when 8032 => read_data_o <= x"0000";
when 8033 => read_data_o <= x"0000";
when 8034 => read_data_o <= x"0000";
when 8035 => read_data_o <= x"0000";
when 8036 => read_data_o <= x"0000";
when 8037 => read_data_o <= x"0000";
when 8038 => read_data_o <= x"0000";
when 8039 => read_data_o <= x"0000";
when 8040 => read_data_o <= x"0000";
when 8041 => read_data_o <= x"0000";
when 8042 => read_data_o <= x"0000";
when 8043 => read_data_o <= x"0000";
when 8044 => read_data_o <= x"0000";
when 8045 => read_data_o <= x"0000";
when 8046 => read_data_o <= x"0000";
when 8047 => read_data_o <= x"0000";
when 8048 => read_data_o <= x"0000";
when 8049 => read_data_o <= x"0000";
when 8050 => read_data_o <= x"0000";
when 8051 => read_data_o <= x"0000";
when 8052 => read_data_o <= x"d770";
when 8053 => read_data_o <= x"041a";
when 8054 => read_data_o <= x"0000";
when 8055 => read_data_o <= x"0000";
when 8056 => read_data_o <= x"002a";
when 8057 => read_data_o <= x"0000";
when 8058 => read_data_o <= x"0000";
when 8059 => read_data_o <= x"0000";
when 8060 => read_data_o <= x"0000";
when 8061 => read_data_o <= x"0000";
when 8062 => read_data_o <= x"a600";
when 8063 => read_data_o <= x"64d5";
when 8064 => read_data_o <= x"0000";
when 8065 => read_data_o <= x"0000";
when 8066 => read_data_o <= x"0000";
when 8067 => read_data_o <= x"0000";
when 8068 => read_data_o <= x"0000";
when 8069 => read_data_o <= x"0000";
when 8070 => read_data_o <= x"0000";
when 8071 => read_data_o <= x"0000";
when 8072 => read_data_o <= x"0000";
when 8073 => read_data_o <= x"0000";
when 8074 => read_data_o <= x"0000";
when 8075 => read_data_o <= x"0000";
when 8076 => read_data_o <= x"0000";
when 8077 => read_data_o <= x"0000";
when 8078 => read_data_o <= x"0000";
when 8079 => read_data_o <= x"0000";
when 8080 => read_data_o <= x"0000";
when 8081 => read_data_o <= x"0000";
when 8082 => read_data_o <= x"0000";
when 8083 => read_data_o <= x"0000";
when 8084 => read_data_o <= x"0000";
when 8085 => read_data_o <= x"0000";
when 8086 => read_data_o <= x"0000";
when 8087 => read_data_o <= x"0000";
when 8088 => read_data_o <= x"0000";
when 8089 => read_data_o <= x"0000";
when 8090 => read_data_o <= x"0000";
when 8091 => read_data_o <= x"0000";
when 8092 => read_data_o <= x"0000";
when 8093 => read_data_o <= x"0000";
when 8094 => read_data_o <= x"0000";
when 8095 => read_data_o <= x"0000";
when 8096 => read_data_o <= x"0000";
when 8097 => read_data_o <= x"0000";
when 8098 => read_data_o <= x"0000";
when 8099 => read_data_o <= x"0000";
when 8100 => read_data_o <= x"0000";
when 8101 => read_data_o <= x"0000";
when 8102 => read_data_o <= x"0000";
when 8103 => read_data_o <= x"0000";
when 8104 => read_data_o <= x"0000";
when 8105 => read_data_o <= x"0000";
when 8106 => read_data_o <= x"0000";
when 8107 => read_data_o <= x"0000";
when 8108 => read_data_o <= x"0000";
when 8109 => read_data_o <= x"0000";
when 8110 => read_data_o <= x"0000";
when 8111 => read_data_o <= x"0000";
when 8112 => read_data_o <= x"0000";
when 8113 => read_data_o <= x"0000";
when 8114 => read_data_o <= x"0000";
when 8115 => read_data_o <= x"0000";
when 8116 => read_data_o <= x"0000";
when 8117 => read_data_o <= x"0000";
when 8118 => read_data_o <= x"0000";
when 8119 => read_data_o <= x"0000";
when 8120 => read_data_o <= x"0000";
when 8121 => read_data_o <= x"0000";
when 8122 => read_data_o <= x"0000";
when 8123 => read_data_o <= x"0000";
when 8124 => read_data_o <= x"0000";
when 8125 => read_data_o <= x"0000";
when 8126 => read_data_o <= x"0000";
when 8127 => read_data_o <= x"0000";
when 8128 => read_data_o <= x"0000";
when 8129 => read_data_o <= x"0000";
when 8130 => read_data_o <= x"7069";
when 8131 => read_data_o <= x"0078";
when 8132 => read_data_o <= x"d770";
when 8133 => read_data_o <= x"041a";
when 8134 => read_data_o <= x"0000";
when 8135 => read_data_o <= x"0000";
when 8136 => read_data_o <= x"002b";
when 8137 => read_data_o <= x"0000";
when 8138 => read_data_o <= x"0000";
when 8139 => read_data_o <= x"0000";
when 8140 => read_data_o <= x"0000";
when 8141 => read_data_o <= x"0000";
when 8142 => read_data_o <= x"0000";
when 8143 => read_data_o <= x"0000";
when 8144 => read_data_o <= x"0000";
when 8145 => read_data_o <= x"0000";
when 8146 => read_data_o <= x"0000";
when 8147 => read_data_o <= x"0000";
when 8148 => read_data_o <= x"0000";
when 8149 => read_data_o <= x"0000";
when 8150 => read_data_o <= x"0000";
when 8151 => read_data_o <= x"0000";
when 8152 => read_data_o <= x"0000";
when 8153 => read_data_o <= x"0000";
when 8154 => read_data_o <= x"0000";
when 8155 => read_data_o <= x"0000";
when 8156 => read_data_o <= x"0000";
when 8157 => read_data_o <= x"0000";
when 8158 => read_data_o <= x"0000";
when 8159 => read_data_o <= x"0000";
when 8160 => read_data_o <= x"0000";
when 8161 => read_data_o <= x"0000";
when 8162 => read_data_o <= x"0000";
when 8163 => read_data_o <= x"0000";
when 8164 => read_data_o <= x"0000";
when 8165 => read_data_o <= x"0000";
when 8166 => read_data_o <= x"0000";
when 8167 => read_data_o <= x"0000";
when 8168 => read_data_o <= x"0000";
when 8169 => read_data_o <= x"0000";
when 8170 => read_data_o <= x"0000";
when 8171 => read_data_o <= x"0000";
when 8172 => read_data_o <= x"0000";
when 8173 => read_data_o <= x"0000";
when 8174 => read_data_o <= x"0000";
when 8175 => read_data_o <= x"0000";
when 8176 => read_data_o <= x"0000";
when 8177 => read_data_o <= x"0000";
when 8178 => read_data_o <= x"0000";
when 8179 => read_data_o <= x"0000";
when 8180 => read_data_o <= x"0000";
when 8181 => read_data_o <= x"0000";
when 8182 => read_data_o <= x"0000";
when 8183 => read_data_o <= x"0000";
when 8184 => read_data_o <= x"0000";
when 8185 => read_data_o <= x"0000";
when 8186 => read_data_o <= x"0000";
when 8187 => read_data_o <= x"0000";
when 8188 => read_data_o <= x"0000";
when 8189 => read_data_o <= x"0000";
when 8190 => read_data_o <= x"0000";
when 8191 => read_data_o <= x"0000";

				when others => read_data_o <= x"a000";
			end case;
		end if;
	end process;

end rtl;
