library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library unisim;
use unisim.Vcomponents.all;
library unimacro;
use unimacro.Vcomponents.all;
entity fontrom is port(
	clk_i  : in std_logic;
	addr_i : in integer;
	data_o : out std_logic_vector(0 downto 0));
end fontrom;

architecture rtl of fontrom is

signal rom_addr_s: std_logic_vector(14 downto 0);
signal rom_data_s: std_logic_vector(31 downto 0);
signal data0_s: std_logic_vector(0 downto 0);
signal data1_s: std_logic_vector(0 downto 0);
begin

rom0: RAMB16_S1
	generic map(
		INIT_00 => X"0008006001800600180060000000000000000000000000000000000000000000",
		INIT_01 => X"00000000000000000000000000000000000CC066019800000000180060000002",
		INIT_02 => X"36007E006C199836C07E0060000019806607FE1FF819806607FE1FF819806600",
		INIT_03 => X"000000000000E186CC1B603B001800DC06D83361870000000006007E036C1998",
		INIT_04 => X"00000000000001C00C003800E0000018C036017415D05DC17F08A803E01FC041",
		INIT_05 => X"18003800001C0018003000600180060018006003001801C00000000000000000",
		INIT_06 => X"1DB80F003C076E19980600180000000003801800C00600180060018006000C00",
		INIT_07 => X"000000000000000018006001803FC0FF00600180060000000000000600180666",
		INIT_08 => X"000000FFF3FFC00000000000000000000007003000E000000000000000000000",
		INIT_09 => X"6003000800000000003800E00000000000000000000000000000000000000000",
		INIT_0A => X"01980C3030C0C3030C0C3030C06600F0000C006003001800C006003001800C00",
		INIT_0B => X"006060C301F800000000FF006001800600180060019007801C0060000000003C",
		INIT_0C => X"7E030C18186000C001F00C006060C301F800000001FF80060070070070030018",
		INIT_0D => X"07F800600183FE000000006001801FF8186063019806C01E0070018000000000",
		INIT_0E => X"007E030C18186060C381F6001800C0C601F0000000007E030C18186001800300",
		INIT_0F => X"F80C306060C301F80000000006001800C006003001800C0060018007FE000000",
		INIT_10 => X"00003E018C0C006001BE070C18186060C301F8000000007E030C18186060C301",
		INIT_11 => X"00E000000000000000000000003800E0000000003800E0000000000000000000",
		INIT_12 => X"00080030006000C0018006003001800C00200000000007003000E00000000038",
		INIT_13 => X"6000C001800300040000000000000003FC0FF000000003FC0FF0000000000000",
		INIT_14 => X"000000003800E000000E0030038018006060C301F8000001000C006003001800",
		INIT_15 => X"C0C3030C066019803C00F0000019802C02F40BD03FC066006003C00F00180000",
		INIT_16 => X"F0000000007F830618186060C181FE0C186060C181FE0000000181860618183F",
		INIT_17 => X"6061818606181830606180FE000000007C031818300060018006001860C0C601",
		INIT_18 => X"87FE00000001FF8006001800600181FE001800600187FE000000003F81860C18",
		INIT_19 => X"306061F18006001860C0C601F000000000018006001800607F80060018006001",
		INIT_1A => X"1801F800000001818606181860618187FE1818606181860600000001BC071818",
		INIT_1B => X"0C006001800600180060018007F0000000007E00600180060018006001800600",
		INIT_1C => X"60018006000000018186060C18186031807E03181860C18606000000003F0186",
		INIT_1D => X"06181860619986F61E7870E181840200000001FF800600180060018006001800",
		INIT_1E => X"30C06600F0000000018186061C187861B1866618D861E1838606000000018186",
		INIT_1F => X"8006001800607F830618186060C181FE000000003C01980C3060618186061818",
		INIT_20 => X"186060C181FE0C0038003C01D80DB06061818606181830C06600F00000000001",
		INIT_21 => X"7E030C18186000C001F800300060C301F8000000018186060C1818607F830618",
		INIT_22 => X"181860618186060000000018006001800600180060018006001807FE00000000",
		INIT_23 => X"003C00F006601980C3030C0C306061818606000000003C01980C306061818606",
		INIT_24 => X"6003C01980C30606000000006601980FF036C0DB066619986061818606000000",
		INIT_25 => X"0000180060018006001800F0066030C1818606000000018186060C3019803C00",
		INIT_26 => X"0018006001800601F800000001FF800C006003001800C0060030018007FE0000",
		INIT_27 => X"006000C00180030006000C00180030006000C00100001F800600180060018006",
		INIT_28 => X"00030C06600F0018000000001F8060018006001800600180060018006001F830",
		INIT_29 => X"1FF87FE000000000000000000000000000000000000000000000000000000000",
		INIT_2A => X"C1FE06000C101FC00000000000000000000000000000000000038003001C0070",
		INIT_2B => X"00000000003D830E1818606181860E0CD81E6001800600000001BE078C1C1860",
		INIT_2C => X"60618186061C306F01800600000000003C030C081800600182060C300F000000",
		INIT_2D => X"078000000000FC060C00180061FF860618301F00000000000000019E06CC1C18",
		INIT_2E => X"3070618186061C306F0000000000000000180060018006001803F80180060030",
		INIT_2F => X"180060000000018186061818606181860E0CD81E6001800607F030618006781B",
		INIT_30 => X"0180060018006001F00000180060000000001800600180060018006001F00000",
		INIT_31 => X"0018007C00000001818386039803E03983861818006001800600780300180060",
		INIT_32 => X"66199866619986661BB83BA00000000000000018006001800600180060018006",
		INIT_33 => X"0F00000000000000018186061818606181860E0CD81E60000000000000019986",
		INIT_34 => X"830E1818606181860E0CD81E60000000000000003C030C181860618186060C30",
		INIT_35 => X"D83E60000000180060019E06CC1C1860618186061C306F00000000001800603D",
		INIT_36 => X"7F060618003C000F00060C181FC0000000000000000180060018006001860E18",
		INIT_37 => X"1818606000000000000001E000C00180060018006001803F8018004000000000",
		INIT_38 => X"001800F006601980C3030C18186060000000000000019E06CC1C186061818606",
		INIT_39 => X"980C306060000000000000006601980FF036C199866618186060000000000000",
		INIT_3A => X"30618006781B307061818606181860600000000000000181830C06600F003C01",
		INIT_3B => X"013213B0220034018C00000001FF001800C006003001800C007FC000000007F0",
		INIT_3C => X"800600180060018006001800600180060018006000001F80FF0606118836C018",
		INIT_3D => X"0000000F106EC11E000030188F30E6040E0700B0119E00CD1818B3006844CC01",
		INIT_3E => X"004844404B80F60DF85EE0F18FEE0FF80D400E00000000000000000000000000",
		INIT_3F => X"404101040220070000000000000F007E01E807200F001800F001800600000000")
	port map(
		SSR => '0',
		DI => "0",
		EN => '1',
		WE => '0',
		CLK => clk_i,
		ADDR => rom_addr_s(13 downto 0),
		DO => data0_s
	);

rom1: RAMB16_S1
	generic map(
		INIT_00 => X"0000001F8018006007E03FC08102F400000000000000000007003E0070022010",
		INIT_01 => X"6F217883DE007800C0030000000036C1E7836C03C036C06600C0000000000000",
		INIT_02 => X"000000000F807F018C0C183160C9838E07F01FC03E000000001F80C2052E1428",
		INIT_03 => X"645FF0DB46DA06D00000000000000021008201B003004F217302E00240090018",
		INIT_04 => X"000000000000800700F801800F006003000800600100000000001FF0BB45ED0A",
		INIT_05 => X"17C859E1EB06BC0CE00F800C00000000000008005002E017C03E000000000000",
		INIT_06 => X"D3FFCFFF00005002A00540050008005D80C900D8000000000000001C008C02CC",
		INIT_07 => X"0000000600180000000000000000003FFC801200C9FD242C90D242C90D27ECBF",
		INIT_08 => X"00000000000000000003001C00A007002801400E001000000000000000000000",
		INIT_09 => X"86A619582AA11500A219186A619586AE0000000000007002600B803E00700000",
		INIT_0A => X"FC3572A9C1FC00005552AA85552AA8555238CBEF0E38555071C71C11502A2191",
		INIT_0B => X"AA85552AA800015542AB2FFC3572A9C1FC11502A219186061AB800015542AB2F",
		INIT_0C => X"003800A001800000000000000000000000000000000FF05561FF800000005552",
		INIT_0D => X"01FF87B413F85FE17F87B41FF83FC00000000000006003800A003800A003800A",
		INIT_0E => X"EA1554AAA1554AAA0444444044444405C4494064446404444440444444000000",
		INIT_0F => X"04001B013C07E007C07D83D00F6018000000001554AAA1554AAA15D4A9A1654A",
		INIT_10 => X"07C01F000001C00700000008006003F01F601BC07F01A4038007000000000000",
		INIT_11 => X"0000000000F8063010406300F800000000000000000057C0BF05000FC05F0080",
		INIT_12 => X"FF00000FF06F60FF00000E7073819C84E6073839C00E0072001800E000000000",
		INIT_13 => X"00000F807F018C0C183DE0C183DE04101DC03E00000FF06F60FF00000FF06F60",
		INIT_14 => X"008087271FFC252000000000001F0086007003004C513C86761F6839C0420000",
		INIT_15 => X"38044015405501FC17F03F800E80BA01B001000E001000000000000000000000",
		INIT_16 => X"17A052814A07380FC02B00780E00618366CDFF1FAC3D607B0039019807C01D00",
		INIT_17 => X"0040000073813B06E41EE033007F03B21CC86740E6000007780DC016015A05E8",
		INIT_18 => X"CCCF33FFC7FE02401F805A00F000001B006C01500BA03F8028011007C00E0010",
		INIT_19 => X"3E00001554BEA1C14E021814E021804E021804B021414AAA1EF01B01AD86F633",
		INIT_1A => X"13F07B011E04FC11A007800C000000000F8077018C0F7838E0E383DE06301DC0",
		INIT_1B => X"801E0000070013805801C007481E403E00E000B007C01A003804603BE1FC8278",
		INIT_1C => X"FC0F7003C00F0024006003C006000007700D8036815A05E81FE03F007805400F",
		INIT_1D => X"07000000001EF00F01BD86F612486FE1FF008807F01240FF8070020030018E07",
		INIT_1E => X"83F70FDC11F03BC1F50B6024807C00000000780160073C0D581AA05581AC03E0",
		INIT_1F => X"E863E0070000000007007E03BA09F8D7C1CA036C09B005400E0000182033004C",
		INIT_20 => X"EC01A00F607541BB071C0C703F805701F000000E007C03B81CE0675198836E0D",
		INIT_21 => X"045055206C00E0031C0EE01B006D01BC37D1D54D5717FC15503F807C04601980",
		INIT_22 => X"631C81FA05EC1BB05D80C803200E401F00000C603B00FC03FE0FC83FA0FF03FE",
		INIT_23 => X"EE07F00D401E00000DB03FC08101DC07702040AD03BC00103FC0DB000007807B",
		INIT_24 => X"31C04201D011C46730FF81DC0080070008000000003DE03606FB1BEC4C91AEC3",
		INIT_25 => X"C7771554777088800000000000C3056A0AD011814A851A14A81F800000000000",
		INIT_26 => X"001FF0BB45ED0A645FF09985FF0DB46DA06D000000002221DDC5551DDC7771DD",
		INIT_27 => X"0000000000000000000000000D806301DC0E383760DD838E077018C036000000",
		INIT_28 => X"000005002B015E09E817E0BD81E407F00F0000000000007FE08302541EB83FC0",
		INIT_29 => X"E0F301FA0BF006000000000000158054855E0B700E00DD038800000000000000",
		INIT_2A => X"0000001E00C4062018007901FE03F000D802C00C0000001010011A80F00BF07C",
		INIT_2B => X"1BA06A81BA07180FC01E000000000300CB02280BA03FB07DC60E306801200000",
		INIT_2C => X"C00000001CE0C606F71FBC3FF0FD441B10444000C00000000000000000780310",
		INIT_2D => X"D01DC01400A803E0070008000003600F609783AC05C00F802A00A807F038E1C1",
		INIT_2E => X"00000000000D801403F411D00F805C01F802A0000000000000000D8036007005",
		INIT_2F => X"05D01FC036007002A00F8022000000000F007F03FE1DB87261FF837E03B00600",
		INIT_30 => X"001C000000002E609B027408E82EE0EE027C14E0210004000000000D80140174",
		INIT_31 => X"D402D83EE0F587DC0070038006000000001DC03600D80BE837607F00F801C007",
		INIT_32 => X"0FC03501FE00006300D803E00F801E008C05DA0AB01CC006003000007F00FA01",
		INIT_33 => X"C3EB1FAC7EE0FA8BF0170000000000000000000004001000C003000E007801E0",
		INIT_34 => X"80000000000000001800CC06A61BFC7FE1FA83DE00480000000000006031A0DD",
		INIT_35 => X"FE01500000000000000000000000000000000008819281DE19F01F80F9019000",
		INIT_36 => X"09C81E400000000000110055015407F05FC0FE003600F803C00600003FF864C0",
		INIT_37 => X"007803F01DE067803F00B401E007800C0000000013C09C82D80EB037606B80DA",
		INIT_38 => X"F807E036C0180000000000803B00B80BF817A1BF83E01E607600000000000000",
		INIT_39 => X"18C07E00F30DFC3561E8067A0D780EC01000000000000018036C07E01F81FF81",
		INIT_3A => X"83FE07F00F8000000000000F807F01240E383DE0F7830606301DC03E00000F78",
		INIT_3B => X"000F807301940E183CE0FF83CE07F01CC03E000000006D30DD83FE0D28252094",
		INIT_3C => X"02801C01BC1A418A88D101E01FE0C0C203081C11E27E0E40008003001C03C000",
		INIT_3D => X"00000000000000000000000000000000000000000000040020008004001400A0",
		INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
	port map(
		SSR => '0',
		DI => "0",
		EN => '1',
		WE => '0',
		CLK => clk_i,
		ADDR => rom_addr_s(13 downto 0),
		DO => data1_s);

rom_addr_s <= std_logic_vector(to_unsigned(addr_i, rom_addr_s'length));
data_o <= data1_s when rom_addr_s(14) = '1' else data0_s;
end rtl;
