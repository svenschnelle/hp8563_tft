library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library unisim;
use unisim.Vcomponents.all;
library unimacro;
use unimacro.Vcomponents.all;
entity fontrom is port(
	clk_i  : in std_logic;
	addr_i : in integer;
	data_o : out std_logic_vector(0 downto 0));
end fontrom;

architecture rtl of fontrom is

signal rom_addr_s: std_logic_vector(14 downto 0);
signal rom_data_s: std_logic_vector(31 downto 0);
signal data0_s: std_logic_vector(0 downto 0);
signal data1_s: std_logic_vector(0 downto 0);
begin

rom0: RAMB16_S1
	generic map(
INIT_00 => X"0008006001800600180060000000000000000000000000000000000000000000",
INIT_01 => X"00000000000000000000000000000000000CC066019800000000180060000002",
INIT_02 => X"36007E006C199836C07E0060000019806607FE1FF819806607FE1FF819806600",
INIT_03 => X"000000000000E186CC1B603B001800DC06D83361870000000006007E036C1998",
INIT_04 => X"00000000000001C00C003800E0000018C036017415D05DC17F08A803E01FC041",
INIT_05 => X"18003800001C0018003000600180060018006003001801C00000000000000000",
INIT_06 => X"1DB80F003C076E19980600180000000003801800C00600180060018006000C00",
INIT_07 => X"000000000000000018006001803FC0FF00600180060000000000000600180666",
INIT_08 => X"000000FFF3FFC00000000000000000000007003000E000000000000000000000",
INIT_09 => X"6003000800000000003800E00000000000000000000000000000000000000000",
INIT_0A => X"01980C3030C0C3030C0C3030C06600F0000C006003001800C006003001800C00",
INIT_0B => X"006060C301F800000000FF006001800600180060019007801C0060000000003C",
INIT_0C => X"7E030C18186000C001F00C006060C301F800000001FF80060070070070030018",
INIT_0D => X"07F800600183FE000000006001801FF8186063019806C01E0070018000000000",
INIT_0E => X"007E030C18186060C381F6001800C0C601F0000000007E030C18186001800300",
INIT_0F => X"F80C306060C301F80000000006001800C006003001800C0060018007FE000000",
INIT_10 => X"00003E018C0C006001BE070C18186060C301F8000000007E030C18186060C301",
INIT_11 => X"00E000000000000000000000003800E0000000003800E0000000000000000000",
INIT_12 => X"00080030006000C0018006003001800C00200000000007003000E00000000038",
INIT_13 => X"6000C001800300040000000000000003FC0FF000000003FC0FF0000000000000",
INIT_14 => X"000000003800E000000E0030038018006060C301F8000001000C006003001800",
INIT_15 => X"C0C3030C066019803C00F0000019802C02F40BD03FC066006003C00F00180000",
INIT_16 => X"F0000000007F830618186060C181FE0C186060C181FE0000000181860618183F",
INIT_17 => X"6061818606181830606180FE000000007C031818300060018006001860C0C601",
INIT_18 => X"87FE00000001FF8006001800600181FE001800600187FE000000003F81860C18",
INIT_19 => X"306061F18006001860C0C601F000000000018006001800607F80060018006001",
INIT_1A => X"1801F800000001818606181860618187FE1818606181860600000001BC071818",
INIT_1B => X"0C006001800600180060018007F0000000007E00600180060018006001800600",
INIT_1C => X"60018006000000018186060C18186031807E03181860C18606000000003F0186",
INIT_1D => X"06181860619986F61E7870E181840200000001FF800600180060018006001800",
INIT_1E => X"30C06600F0000000018186061C187861B1866618D861E1838606000000018186",
INIT_1F => X"8006001800607F830618186060C181FE000000003C01980C3060618186061818",
INIT_20 => X"186060C181FE0C0038003C01D80DB06061818606181830C06600F00000000001",
INIT_21 => X"7E030C18186000C001F800300060C301F8000000018186060C1818607F830618",
INIT_22 => X"181860618186060000000018006001800600180060018006001807FE00000000",
INIT_23 => X"003C00F006601980C3030C0C306061818606000000003C01980C306061818606",
INIT_24 => X"6003C01980C30606000000006601980FF036C0DB066619986061818606000000",
INIT_25 => X"0000180060018006001800F0066030C1818606000000018186060C3019803C00",
INIT_26 => X"0018006001800601F800000001FF800C006003001800C0060030018007FE0000",
INIT_27 => X"006000C00180030006000C00180030006000C00100001F800600180060018006",
INIT_28 => X"00030C06600F0018000000001F8060018006001800600180060018006001F830",
INIT_29 => X"1FF87FE000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"C1FE06000C101FC00000000000000000000000000000000000038003001C0070",
INIT_2B => X"00000000003D830E1818606181860E0CD81E6001800600000001BE078C1C1860",
INIT_2C => X"60618186061C306F01800600000000003C030C081800600182060C300F000000",
INIT_2D => X"078000000000FC060C00180061FF860618301F00000000000000019E06CC1C18",
INIT_2E => X"3070618186061C306F0000000000000000180060018006001803F80180060030",
INIT_2F => X"180060000000018186061818606181860E0CD81E6001800607F030618006781B",
INIT_30 => X"0180060018006001F00000180060000000001800600180060018006001F00000",
INIT_31 => X"0018007C00000001818386039803E03983861818006001800600780300180060",
INIT_32 => X"66199866619986661BB83BA00000000000000018006001800600180060018006",
INIT_33 => X"0F00000000000000018186061818606181860E0CD81E60000000000000019986",
INIT_34 => X"830E1818606181860E0CD81E60000000000000003C030C181860618186060C30",
INIT_35 => X"D83E60000000180060019E06CC1C1860618186061C306F00000000001800603D",
INIT_36 => X"7F060618003C000F00060C181FC0000000000000000180060018006001860E18",
INIT_37 => X"1818606000000000000001E000C00180060018006001803F8018004000000000",
INIT_38 => X"001800F006601980C3030C18186060000000000000019E06CC1C186061818606",
INIT_39 => X"980C306060000000000000006601980FF036C199866618186060000000000000",
INIT_3A => X"30618006781B307061818606181860600000000000000181830C06600F003C01",
INIT_3B => X"013213B0220034018C00000001FF001800C006003001800C007FC000000007F0",
INIT_3C => X"800600180060018006001800600180060018006000001F80FF0606118836C018",
INIT_3D => X"0000000F106EC11E000030188F30E6040E0700B0119E00CD1818B3006844CC01",
INIT_3E => X"004844404B80F60DF85EE0F18FEE0FF80D400E00000000000000000000000000",
INIT_3F => X"404101040220070000000000000F007E01E807200F001800F001800600000000")
		port map(
		SSR => '0',
		DI => "0",
		EN => '1',
		WE => '0',
		CLK => clk_i,
		ADDR => rom_addr_s(13 downto 0),
		DO => data0_s
	);

rom1: RAMB16_S1
	generic map(
		INIT_00 => X"0804400E007C00E00000000000000000002F408103FC07E006001801F8000000",
		INIT_01 => X"000000000000030066036C03C036C1E7836C00000000C003001E007BC11E84F6",
		INIT_02 => X"142874A04301F8000000007C03F80FE071C193068C18303180FE01F000000000",
		INIT_03 => X"18009002400740CE84F200C00D80410084000000000000000B605B62DB0FFA26",
		INIT_04 => X"50B7A2DD0FF800000000008006001000C00600F001801F00E001000000000000",
		INIT_05 => X"0000000000007C03E807400A00100000000000003001F007303D60D7879A13E8",
		INIT_06 => X"3340310038000000000000001B009301BA001000A002A005400A0000FFF3FFCB",
		INIT_07 => X"FD37E4B093424B093424BF930048013FFC000000000000000000180060000000",
		INIT_08 => X"0000000000000000000008007002801400E005003800C0000000000000000000",
		INIT_09 => X"00000E007C01D006400E0000000000007561A9865618984500A885541A986561",
		INIT_0A => X"8984540A8838E38E0AAA1C70F7D31C4AAA1554AAA1554AAA00003F83954EAC3F",
		INIT_0B => X"F4D542AA80001D5860618984540A883F83954EAC3FF4D542AA80001554AAA155",
		INIT_0C => X"4AAA00000001FF86AA0FF0000000000000000000000000000000018005001C00",
		INIT_0D => X"5001C005001C005001C00600000000000003FC1FF82DE1FE87FA1FC82DE1FF80",
		INIT_0E => X"00000022222202222220262226029223A0222222022222205552AA85552AA857",
		INIT_0F => X"52A685952BA85552AA85552AA8000000001806F00BC1BE03E007E03C80D80020",
		INIT_10 => X"000000000000E001C02580FE03D806F80FC0060010000000E003800000F803E0",
		INIT_11 => X"0100FA03F000A0FD03EA0000000000000000001F00C602080C601F0000000000",
		INIT_12 => X"00000000070018004E0070039C1CE067213981CE0E700000FF06F60FF00000FF",
		INIT_13 => X"06F60FF00000FF06F60FF000007C03B808207BC18307BC18303180FE01F00000",
		INIT_14 => X"000042039C16F86E613C8A3200C00E006100F8000000000004A43FF8E4E10100",
		INIT_15 => X"0000000000000000000008007000800D805D017001FC0FE83F80AA02A802201C",
		INIT_16 => X"00B803E019809C00DE06BC35F8FFB366C18600701E00D403F01CE052814A05E8",
		INIT_17 => X"17A05A806803B01EE000006702E613384DC0FE00CC07782760DC81CE00000200",
		INIT_18 => X"08007003E008801401FC05D00A803600D800000F005A01F802407FE3FFCCF333",
		INIT_19 => X"CC6F61B580D80F78555282840D201840720184072818407283857D2AA800007C",
		INIT_1A => X"03B80C607BC1C7071C1EF03180EE01F0000000003001E005883F207880DE0FC8",
		INIT_1B => X"1E413F87DC06201C005803E00D0007007C027812E003801A01C800E000007801",
		INIT_1C => X"F002A01E00FC07F817A05A816C01B00EE000006003C006002400F003C00EF03F",
		INIT_1D => X"E071800C00400E01FF02480FE01100FF87F612486F61BD80F00F7800000000E0",
		INIT_1E => X"07C03581AA05581AB03CE006801E000000003E012406D0AF83DC0F883BF0EFC1",
		INIT_1F => X"3200CC041800007002A00D9036C05383EB1F905DC07E00E000000000E007C617",
		INIT_20 => X"B076C1198AE607381DC03E007000000F80EA01FC0E3038E0DD82AE06F0058037",
		INIT_21 => X"019806203E01FC0AA83FE8EAB2AB8BEC3D80B600D8077038C007003604AA0A20",
		INIT_22 => X"7FC0FF05FC13F07FC03F00DC06300000F8027004C01301BA0DD837A05F8138C6",
		INIT_23 => X"DE01E00000DB03FC08003DC0B502040EE03B808103FC0DB000007802B00FE077",
		INIT_24 => X"C375893237D8DF606C07BC000000001000E001003B81FF0CE623880B8042038C",
		INIT_25 => X"000000000001F8152858A15281880B5056A0C3000000000001110EEE2AA8EEE3",
		INIT_26 => X"BB8EEE3BB8AAA3BB844400000000B605B62DB0FFA1990FFA2650B7A2DD0FF800",
		INIT_27 => X"0000006C03180EE071C1BB06EC1C703B80C601B0000000000000000000000000",
		INIT_28 => X"03FC1D782A40C107FE000000000000F00FE02781BD07E817907A80D400A00000",
		INIT_29 => X"0000000000000011C0BB00700ED07AA12A01A8000000000000600FD05F80CF07",
		INIT_2A => X"3E0FD00F01588008080000003003401B000FC07F809E00180460230078000000",
		INIT_2B => X"00000480160C7063BE0DFC05D01440D300C0000000007803F018E05D815605D8",
		INIT_2C => X"08C01E00000000000000000300022208D822BF0FFC3DF8EF6063073800000003",
		INIT_2D => X"83871C0FE015005401F003A035C1E906F006C000001000E007C015002803B80B",
		INIT_2E => X"A00E006C01B00000000000000005401F803A01F00B882FC02801B00000000000",
		INIT_2F => X"00600DC07EC1FF864E1DB87FC0FE00F0000000004401F005400E006C03F80BA0",
		INIT_30 => X"2E802801B00000000020008407283E4077077417102E40D90674000000003800",
		INIT_31 => X"E003801F00FE06EC17D01B006C03B8000000006001C00E003BE1AF077C1B402B",
		INIT_32 => X"805F00FE00000C006003380D505BA031007801F007C01B00C600007F80AC03F0",
		INIT_33 => X"07801E007000C0030008002000000000000000000000E80FD15F077E35F8D7C3",
		INIT_34 => X"BB058C0600000000000012007BC15F87FE3FD865603300180000000000000001",
		INIT_35 => X"0009809F01F80F987B81498110000000000000000000000000000000000A807F",
		INIT_36 => X"03261FFC00006003C01F006C007F03FA0FE02A80AA0088000000000002781390",
		INIT_37 => X"5B01D606EC0D701B413903C8000000003001E007802D00FC01E607B80FC01E00",
		INIT_38 => X"000000000000006E067807C1FD85E81FD01D00DC01000000000018036C07E01F",
		INIT_39 => X"81FF81F807E036C0180000000000000803701EB05E601786AC3FB0CF007E0318",
		INIT_3A => X"1EF000007C03B80C6060C1EF07BC1C702480FE01F0000000000001F00FE07FC1",
		INIT_3B => X"2904A414B07FC1BB0CB6000000007C03380FE073C1FF073C18702980CE01F000",
		INIT_3C => X"0003C03800C0010002707E47883810C0430307F807808B115182583D80380140",
		INIT_3D => X"0500280020010004002000000000000000000000000000000000000000000000",
		INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
	port map(
		SSR => '0',
		DI => "0",
		EN => '1',
		WE => '0',
		CLK => clk_i,
		ADDR => rom_addr_s(13 downto 0),
		DO => data1_s);

rom_addr_s <= std_logic_vector(to_unsigned(addr_i, rom_addr_s'length));
data_o <= data1_s when rom_addr_s(14) = '1' else data0_s;
end rtl;
