library ieee;
use ieee.std_logic_1164.all;

entity testrom is
	port(read_clock_i: in std_logic;
	   read_addr_i: in integer range 0 to 8191;
	   read_data_o: out std_logic_vector(15 downto 0)
);
end testrom;
architecture rtl of testrom is
begin
	process (read_clock_i)
	begin
		if (rising_edge(read_clock_i)) then
			case read_addr_i is
				when 16#0000# => read_data_o <= x"a002";
				when 16#0001# => read_data_o <= x"7318";
				when 16#0002# => read_data_o <= x"0264";
				when 16#0003# => read_data_o <= x"4350";
				when 16#0004# => read_data_o <= x"0264";
				when 16#0005# => read_data_o <= x"72c8";
				when 16#0006# => read_data_o <= x"0200";
				when 16#0007# => read_data_o <= x"4310";
				when 16#0008# => read_data_o <= x"0200";
				when 16#0009# => read_data_o <= x"7318";
				when 16#000a# => read_data_o <= x"019c";
				when 16#000b# => read_data_o <= x"4350";
				when 16#000c# => read_data_o <= x"019c";
				when 16#000d# => read_data_o <= x"72c0";
				when 16#000e# => read_data_o <= x"00f0";
				when 16#000f# => read_data_o <= x"72d0";
				when 16#0010# => read_data_o <= x"00f0";
				when 16#0011# => read_data_o <= x"72c0";
				when 16#0012# => read_data_o <= x"008c";
				when 16#0013# => read_data_o <= x"72d0";
				when 16#0014# => read_data_o <= x"008c";
				when 16#0015# => read_data_o <= x"7318";
				when 16#0016# => read_data_o <= x"0070";
				when 16#0017# => read_data_o <= x"4350";
				when 16#0018# => read_data_o <= x"0070";
				when 16#0019# => read_data_o <= x"72c8";
				when 16#001a# => read_data_o <= x"02e2";
				when 16#001b# => read_data_o <= x"72c8";
				when 16#001c# => read_data_o <= x"02e2";
				when 16#001d# => read_data_o <= x"4350";
				when 16#001e# => read_data_o <= x"02e2";
				when 16#001f# => read_data_o <= x"7350";
				when 16#0020# => read_data_o <= x"02e2";
				when 16#0021# => read_data_o <= x"5350";
				when 16#0022# => read_data_o <= x"02be";
				when 16#0023# => read_data_o <= x"7350";
				when 16#0024# => read_data_o <= x"02be";
				when 16#0025# => read_data_o <= x"42c8";
				when 16#0026# => read_data_o <= x"02be";
				when 16#0027# => read_data_o <= x"72c8";
				when 16#0028# => read_data_o <= x"02be";
				when 16#0029# => read_data_o <= x"52c8";
				when 16#002a# => read_data_o <= x"02e2";
				when 16#002b# => read_data_o <= x"72c8";
				when 16#002c# => read_data_o <= x"02e2";
				when 16#002d# => read_data_o <= x"72c8";
				when 16#002e# => read_data_o <= x"02e2";
				when 16#002f# => read_data_o <= x"4350";
				when 16#0030# => read_data_o <= x"02e2";
				when 16#0031# => read_data_o <= x"7350";
				when 16#0032# => read_data_o <= x"02e2";
				when 16#0033# => read_data_o <= x"5350";
				when 16#0034# => read_data_o <= x"02be";
				when 16#0035# => read_data_o <= x"7350";
				when 16#0036# => read_data_o <= x"02be";
				when 16#0037# => read_data_o <= x"42c8";
				when 16#0038# => read_data_o <= x"02be";
				when 16#0039# => read_data_o <= x"72c8";
				when 16#003a# => read_data_o <= x"02be";
				when 16#003b# => read_data_o <= x"52c8";
				when 16#003c# => read_data_o <= x"02e2";
				when 16#003d# => read_data_o <= x"62c0";
				when 16#003e# => read_data_o <= x"0294";
				when 16#003f# => read_data_o <= x"c1e5";
				when 16#0040# => read_data_o <= x"c204";
				when 16#0041# => read_data_o <= x"c1c5";
				when 16#0042# => read_data_o <= x"c02b";
				when 16#0043# => read_data_o <= x"c1ef";
				when 16#0044# => read_data_o <= x"c189";
				when 16#0045# => read_data_o <= x"c1a8";
				when 16#0046# => read_data_o <= x"c160";
				when 16#0047# => read_data_o <= x"62c0";
				when 16#0048# => read_data_o <= x"027c";
				when 16#0049# => read_data_o <= x"c137";
				when 16#004a# => read_data_o <= x"c1f6";
				when 16#004b# => read_data_o <= x"c1ef";
				when 16#004c# => read_data_o <= x"c1ba";
				when 16#004d# => read_data_o <= x"c02b";
				when 16#004e# => read_data_o <= x"c1a8";
				when 16#004f# => read_data_o <= x"c137";
				when 16#0050# => read_data_o <= x"c1b2";
				when 16#0051# => read_data_o <= x"a0ca";
				when 16#0052# => read_data_o <= x"0000";
				when 16#0053# => read_data_o <= x"0000";
				when 16#0054# => read_data_o <= x"0000";
				when 16#0055# => read_data_o <= x"0000";
				when 16#0056# => read_data_o <= x"0000";
				when 16#0057# => read_data_o <= x"0000";
				when 16#0058# => read_data_o <= x"0000";
				when 16#0059# => read_data_o <= x"0000";
				when 16#005a# => read_data_o <= x"0000";
				when 16#005b# => read_data_o <= x"0000";
				when 16#005c# => read_data_o <= x"0000";
				when 16#005d# => read_data_o <= x"0000";
				when 16#005e# => read_data_o <= x"0000";
				when 16#005f# => read_data_o <= x"0000";
				when 16#0060# => read_data_o <= x"0000";
				when 16#0061# => read_data_o <= x"0000";
				when 16#0062# => read_data_o <= x"0000";
				when 16#0063# => read_data_o <= x"0000";
				when 16#0064# => read_data_o <= x"0000";
				when 16#0065# => read_data_o <= x"0094";
				when 16#0066# => read_data_o <= x"02dc";
				when 16#0067# => read_data_o <= x"d02b";
				when 16#0068# => read_data_o <= x"d02b";
				when 16#0069# => read_data_o <= x"d1e5";
				when 16#006a# => read_data_o <= x"d204";
				when 16#006b# => read_data_o <= x"d160";
				when 16#006c# => read_data_o <= x"d160";
				when 16#006d# => read_data_o <= x"d1c5";
				when 16#006e# => read_data_o <= x"d02b";
				when 16#006f# => read_data_o <= x"72c0";
				when 16#0070# => read_data_o <= x"0294";
				when 16#0071# => read_data_o <= x"d1e5";
				when 16#0072# => read_data_o <= x"d204";
				when 16#0073# => read_data_o <= x"d1c5";
				when 16#0074# => read_data_o <= x"d02b";
				when 16#0075# => read_data_o <= x"d1ef";
				when 16#0076# => read_data_o <= x"d189";
				when 16#0077# => read_data_o <= x"d1a8";
				when 16#0078# => read_data_o <= x"d160";
				when 16#0079# => read_data_o <= x"72c0";
				when 16#007a# => read_data_o <= x"027c";
				when 16#007b# => read_data_o <= x"d137";
				when 16#007c# => read_data_o <= x"d1f6";
				when 16#007d# => read_data_o <= x"d1ef";
				when 16#007e# => read_data_o <= x"d1ba";
				when 16#007f# => read_data_o <= x"d02b";
				when 16#0080# => read_data_o <= x"d1a8";
				when 16#0081# => read_data_o <= x"d137";
				when 16#0082# => read_data_o <= x"d1b2";
				when 16#0083# => read_data_o <= x"72c0";
				when 16#0084# => read_data_o <= x"0230";
				when 16#0085# => read_data_o <= x"d02b";
				when 16#0086# => read_data_o <= x"d02b";
				when 16#0087# => read_data_o <= x"d02b";
				when 16#0088# => read_data_o <= x"d1e5";
				when 16#0089# => read_data_o <= x"d204";
				when 16#008a# => read_data_o <= x"d160";
				when 16#008b# => read_data_o <= x"d160";
				when 16#008c# => read_data_o <= x"d1c5";
				when 16#008d# => read_data_o <= x"72c0";
				when 16#008e# => read_data_o <= x"0218";
				when 16#008f# => read_data_o <= x"d14e";
				when 16#0090# => read_data_o <= x"d1ba";
				when 16#0091# => read_data_o <= x"d1b2";
				when 16#0092# => read_data_o <= x"d1ef";
				when 16#0093# => read_data_o <= x"d02b";
				when 16#0094# => read_data_o <= x"d1e5";
				when 16#0095# => read_data_o <= x"d174";
				when 16#0096# => read_data_o <= x"d1a2";
				when 16#0097# => read_data_o <= x"72c0";
				when 16#0098# => read_data_o <= x"01cc";
				when 16#0099# => read_data_o <= x"d02b";
				when 16#009a# => read_data_o <= x"d02b";
				when 16#009b# => read_data_o <= x"d02b";
				when 16#009c# => read_data_o <= x"d02b";
				when 16#009d# => read_data_o <= x"d174";
				when 16#009e# => read_data_o <= x"d137";
				when 16#009f# => read_data_o <= x"d1ef";
				when 16#00a0# => read_data_o <= x"d160";
				when 16#00a1# => read_data_o <= x"72c0";
				when 16#00a2# => read_data_o <= x"01b4";
				when 16#00a3# => read_data_o <= x"d02b";
				when 16#00a4# => read_data_o <= x"d02b";
				when 16#00a5# => read_data_o <= x"d1ba";
				when 16#00a6# => read_data_o <= x"d1b2";
				when 16#00a7# => read_data_o <= x"d02b";
				when 16#00a8# => read_data_o <= x"d1ba";
				when 16#00a9# => read_data_o <= x"d16b";
				when 16#00aa# => read_data_o <= x"d16b";
				when 16#00ab# => read_data_o <= x"72c0";
				when 16#00ac# => read_data_o <= x"0168";
				when 16#00ad# => read_data_o <= x"d02b";
				when 16#00ae# => read_data_o <= x"d02b";
				when 16#00af# => read_data_o <= x"d02b";
				when 16#00b0# => read_data_o <= x"d174";
				when 16#00b1# => read_data_o <= x"d137";
				when 16#00b2# => read_data_o <= x"d1ef";
				when 16#00b3# => read_data_o <= x"d160";
				when 16#00b4# => read_data_o <= x"d157";
				when 16#00b5# => read_data_o <= x"72c0";
				when 16#00b6# => read_data_o <= x"0150";
				when 16#00b7# => read_data_o <= x"d02b";
				when 16#00b8# => read_data_o <= x"d02b";
				when 16#00b9# => read_data_o <= x"d02b";
				when 16#00ba# => read_data_o <= x"d1fe";
				when 16#00bb# => read_data_o <= x"d189";
				when 16#00bc# => read_data_o <= x"d157";
				when 16#00bd# => read_data_o <= x"d160";
				when 16#00be# => read_data_o <= x"d1ba";
				when 16#00bf# => read_data_o <= x"72c0";
				when 16#00c0# => read_data_o <= x"0104";
				when 16#00c1# => read_data_o <= x"d02b";
				when 16#00c2# => read_data_o <= x"d157";
				when 16#00c3# => read_data_o <= x"d1a2";
				when 16#00c4# => read_data_o <= x"d215";
				when 16#00c5# => read_data_o <= x"d02b";
				when 16#00c6# => read_data_o <= x"d1e5";
				when 16#00c7# => read_data_o <= x"d204";
				when 16#00c8# => read_data_o <= x"d1c5";
				when 16#00c9# => read_data_o <= x"72c0";
				when 16#00ca# => read_data_o <= x"00ec";
				when 16#00cb# => read_data_o <= x"d225";
				when 16#00cc# => read_data_o <= x"d02b";
				when 16#00cd# => read_data_o <= x"d02b";
				when 16#00ce# => read_data_o <= x"d02b";
				when 16#00cf# => read_data_o <= x"d02b";
				when 16#00d0# => read_data_o <= x"d0a8";
				when 16#00d1# => read_data_o <= x"d2ec";
				when 16#00d2# => read_data_o <= x"d230";
				when 16#00d3# => read_data_o <= x"72c0";
				when 16#00d4# => read_data_o <= x"00a0";
				when 16#00d5# => read_data_o <= x"d02b";
				when 16#00d6# => read_data_o <= x"d157";
				when 16#00d7# => read_data_o <= x"d1a2";
				when 16#00d8# => read_data_o <= x"d215";
				when 16#00d9# => read_data_o <= x"d02b";
				when 16#00da# => read_data_o <= x"d1e5";
				when 16#00db# => read_data_o <= x"d204";
				when 16#00dc# => read_data_o <= x"d1c5";
				when 16#00dd# => read_data_o <= x"72c0";
				when 16#00de# => read_data_o <= x"0088";
				when 16#00df# => read_data_o <= x"d02b";
				when 16#00e0# => read_data_o <= x"d02b";
				when 16#00e1# => read_data_o <= x"d1ba";
				when 16#00e2# => read_data_o <= x"d1b2";
				when 16#00e3# => read_data_o <= x"d02b";
				when 16#00e4# => read_data_o <= x"d1ba";
				when 16#00e5# => read_data_o <= x"d16b";
				when 16#00e6# => read_data_o <= x"d16b";
				when 16#00e7# => read_data_o <= x"a1d0";
				when 16#00e8# => read_data_o <= x"72c0";
				when 16#00e9# => read_data_o <= x"0030";
				when 16#00ea# => read_data_o <= x"d02b";
				when 16#00eb# => read_data_o <= x"d02b";
				when 16#00ec# => read_data_o <= x"d02b";
				when 16#00ed# => read_data_o <= x"d02b";
				when 16#00ee# => read_data_o <= x"d02b";
				when 16#00ef# => read_data_o <= x"d02b";
				when 16#00f0# => read_data_o <= x"d02b";
				when 16#00f1# => read_data_o <= x"d02b";
				when 16#00f2# => read_data_o <= x"72c0";
				when 16#00f3# => read_data_o <= x"0050";
				when 16#00f4# => read_data_o <= x"d02b";
				when 16#00f5# => read_data_o <= x"d02b";
				when 16#00f6# => read_data_o <= x"d02b";
				when 16#00f7# => read_data_o <= x"d02b";
				when 16#00f8# => read_data_o <= x"d02b";
				when 16#00f9# => read_data_o <= x"d02b";
				when 16#00fa# => read_data_o <= x"d02b";
				when 16#00fb# => read_data_o <= x"d02b";
				when 16#00fc# => read_data_o <= x"2403";
				when 16#00fd# => read_data_o <= x"7060";
				when 16#00fe# => read_data_o <= x"01e8";
				when 16#00ff# => read_data_o <= x"d02b";
				when 16#0100# => read_data_o <= x"d02b";
				when 16#0101# => read_data_o <= x"d02b";
				when 16#0102# => read_data_o <= x"d02b";
				when 16#0103# => read_data_o <= x"d02b";
				when 16#0104# => read_data_o <= x"d02b";
				when 16#0105# => read_data_o <= x"d02b";
				when 16#0106# => read_data_o <= x"d02b";
				when 16#0107# => read_data_o <= x"d02b";
				when 16#0108# => read_data_o <= x"d02b";
				when 16#0109# => read_data_o <= x"d02b";
				when 16#010a# => read_data_o <= x"d02b";
				when 16#010b# => read_data_o <= x"d02b";
				when 16#010c# => read_data_o <= x"d02b";
				when 16#010d# => read_data_o <= x"d02b";
				when 16#010e# => read_data_o <= x"d02b";
				when 16#010f# => read_data_o <= x"d02b";
				when 16#0110# => read_data_o <= x"d02b";
				when 16#0111# => read_data_o <= x"d02b";
				when 16#0112# => read_data_o <= x"d02b";
				when 16#0113# => read_data_o <= x"d02b";
				when 16#0114# => read_data_o <= x"d02b";
				when 16#0115# => read_data_o <= x"d02b";
				when 16#0116# => read_data_o <= x"d02b";
				when 16#0117# => read_data_o <= x"d02b";
				when 16#0118# => read_data_o <= x"d02b";
				when 16#0119# => read_data_o <= x"d02b";
				when 16#011a# => read_data_o <= x"d02b";
				when 16#011b# => read_data_o <= x"d02b";
				when 16#011c# => read_data_o <= x"d02b";
				when 16#011d# => read_data_o <= x"d02b";
				when 16#011e# => read_data_o <= x"d02b";
				when 16#011f# => read_data_o <= x"7060";
				when 16#0120# => read_data_o <= x"0202";
				when 16#0121# => read_data_o <= x"d02b";
				when 16#0122# => read_data_o <= x"d02b";
				when 16#0123# => read_data_o <= x"d02b";
				when 16#0124# => read_data_o <= x"d02b";
				when 16#0125# => read_data_o <= x"d02b";
				when 16#0126# => read_data_o <= x"d02b";
				when 16#0127# => read_data_o <= x"d02b";
				when 16#0128# => read_data_o <= x"d02b";
				when 16#0129# => read_data_o <= x"d02b";
				when 16#012a# => read_data_o <= x"d02b";
				when 16#012b# => read_data_o <= x"d02b";
				when 16#012c# => read_data_o <= x"d02b";
				when 16#012d# => read_data_o <= x"d02b";
				when 16#012e# => read_data_o <= x"d02b";
				when 16#012f# => read_data_o <= x"d02b";
				when 16#0130# => read_data_o <= x"d02b";
				when 16#0131# => read_data_o <= x"d02b";
				when 16#0132# => read_data_o <= x"d02b";
				when 16#0133# => read_data_o <= x"d02b";
				when 16#0134# => read_data_o <= x"d02b";
				when 16#0135# => read_data_o <= x"d02b";
				when 16#0136# => read_data_o <= x"d02b";
				when 16#0137# => read_data_o <= x"d02b";
				when 16#0138# => read_data_o <= x"d02b";
				when 16#0139# => read_data_o <= x"d02b";
				when 16#013a# => read_data_o <= x"d02b";
				when 16#013b# => read_data_o <= x"d02b";
				when 16#013c# => read_data_o <= x"d02b";
				when 16#013d# => read_data_o <= x"d02b";
				when 16#013e# => read_data_o <= x"d02b";
				when 16#013f# => read_data_o <= x"d02b";
				when 16#0140# => read_data_o <= x"d02b";
				when 16#0141# => read_data_o <= x"7060";
				when 16#0142# => read_data_o <= x"0224";
				when 16#0143# => read_data_o <= x"d0a8";
				when 16#0144# => read_data_o <= x"d08c";
				when 16#0145# => read_data_o <= x"d095";
				when 16#0146# => read_data_o <= x"d095";
				when 16#0147# => read_data_o <= x"d02b";
				when 16#0148# => read_data_o <= x"d2dc";
				when 16#0149# => read_data_o <= x"d269";
				when 16#014a# => read_data_o <= x"d258";
				when 16#014b# => read_data_o <= x"d02b";
				when 16#014c# => read_data_o <= x"d02b";
				when 16#014d# => read_data_o <= x"d02b";
				when 16#014e# => read_data_o <= x"d02b";
				when 16#014f# => read_data_o <= x"d02b";
				when 16#0150# => read_data_o <= x"d02b";
				when 16#0151# => read_data_o <= x"d02b";
				when 16#0152# => read_data_o <= x"d02b";
				when 16#0153# => read_data_o <= x"d02b";
				when 16#0154# => read_data_o <= x"d02b";
				when 16#0155# => read_data_o <= x"d02b";
				when 16#0156# => read_data_o <= x"7060";
				when 16#0157# => read_data_o <= x"023e";
				when 16#0158# => read_data_o <= x"d1e5";
				when 16#0159# => read_data_o <= x"d204";
				when 16#015a# => read_data_o <= x"d160";
				when 16#015b# => read_data_o <= x"d160";
				when 16#015c# => read_data_o <= x"d1c5";
				when 16#015d# => read_data_o <= x"d1ef";
				when 16#015e# => read_data_o <= x"d189";
				when 16#015f# => read_data_o <= x"d1a8";
				when 16#0160# => read_data_o <= x"d160";
				when 16#0161# => read_data_o <= x"d02b";
				when 16#0162# => read_data_o <= x"d02b";
				when 16#0163# => read_data_o <= x"d02b";
				when 16#0164# => read_data_o <= x"d02b";
				when 16#0165# => read_data_o <= x"d02b";
				when 16#0166# => read_data_o <= x"d02b";
				when 16#0167# => read_data_o <= x"d02b";
				when 16#0168# => read_data_o <= x"d02b";
				when 16#0169# => read_data_o <= x"d02b";
				when 16#016a# => read_data_o <= x"d02b";
				when 16#016b# => read_data_o <= x"71b2";
				when 16#016c# => read_data_o <= x"02ba";
				when 16#016d# => read_data_o <= x"d02b";
				when 16#016e# => read_data_o <= x"d02b";
				when 16#016f# => read_data_o <= x"d02b";
				when 16#0170# => read_data_o <= x"d02b";
				when 16#0171# => read_data_o <= x"d02b";
				when 16#0172# => read_data_o <= x"d02b";
				when 16#0173# => read_data_o <= x"d02b";
				when 16#0174# => read_data_o <= x"d02b";
				when 16#0175# => read_data_o <= x"d02b";
				when 16#0176# => read_data_o <= x"d02b";
				when 16#0177# => read_data_o <= x"d02b";
				when 16#0178# => read_data_o <= x"d02b";
				when 16#0179# => read_data_o <= x"d02b";
				when 16#017a# => read_data_o <= x"d02b";
				when 16#017b# => read_data_o <= x"d02b";
				when 16#017c# => read_data_o <= x"d02b";
				when 16#017d# => read_data_o <= x"71b2";
				when 16#017e# => read_data_o <= x"029c";
				when 16#017f# => read_data_o <= x"d02b";
				when 16#0180# => read_data_o <= x"d02b";
				when 16#0181# => read_data_o <= x"d02b";
				when 16#0182# => read_data_o <= x"d02b";
				when 16#0183# => read_data_o <= x"d02b";
				when 16#0184# => read_data_o <= x"d02b";
				when 16#0185# => read_data_o <= x"d02b";
				when 16#0186# => read_data_o <= x"d02b";
				when 16#0187# => read_data_o <= x"d02b";
				when 16#0188# => read_data_o <= x"d02b";
				when 16#0189# => read_data_o <= x"d02b";
				when 16#018a# => read_data_o <= x"d02b";
				when 16#018b# => read_data_o <= x"d02b";
				when 16#018c# => read_data_o <= x"d02b";
				when 16#018d# => read_data_o <= x"d02b";
				when 16#018e# => read_data_o <= x"d02b";
				when 16#018f# => read_data_o <= x"7040";
				when 16#0190# => read_data_o <= x"0030";
				when 16#0191# => read_data_o <= x"d02b";
				when 16#0192# => read_data_o <= x"d1da";
				when 16#0193# => read_data_o <= x"d140";
				when 16#0194# => read_data_o <= x"d204";
				when 16#0195# => read_data_o <= x"d02b";
				when 16#0196# => read_data_o <= x"d0a1";
				when 16#0197# => read_data_o <= x"d095";
				when 16#0198# => read_data_o <= x"d29c";
				when 16#0199# => read_data_o <= x"d17f";
				when 16#019a# => read_data_o <= x"d30c";
				when 16#019b# => read_data_o <= x"d02b";
				when 16#019c# => read_data_o <= x"7110";
				when 16#019d# => read_data_o <= x"0030";
				when 16#019e# => read_data_o <= x"d02b";
				when 16#019f# => read_data_o <= x"d1fe";
				when 16#01a0# => read_data_o <= x"d140";
				when 16#01a1# => read_data_o <= x"d204";
				when 16#01a2# => read_data_o <= x"d02b";
				when 16#01a3# => read_data_o <= x"d0a1";
				when 16#01a4# => read_data_o <= x"d095";
				when 16#01a5# => read_data_o <= x"d29c";
				when 16#01a6# => read_data_o <= x"d17f";
				when 16#01a7# => read_data_o <= x"d30c";
				when 16#01a8# => read_data_o <= x"d02b";
				when 16#01a9# => read_data_o <= x"71f0";
				when 16#01aa# => read_data_o <= x"0030";
				when 16#01ab# => read_data_o <= x"d074";
				when 16#01ac# => read_data_o <= x"d1e5";
				when 16#01ad# => read_data_o <= x"d204";
				when 16#01ae# => read_data_o <= x"d1c5";
				when 16#01af# => read_data_o <= x"d02b";
				when 16#01b0# => read_data_o <= x"d0a8";
				when 16#01b1# => read_data_o <= x"d08c";
				when 16#01b2# => read_data_o <= x"d095";
				when 16#01b3# => read_data_o <= x"d095";
				when 16#01b4# => read_data_o <= x"d2dc";
				when 16#01b5# => read_data_o <= x"d269";
				when 16#01b6# => read_data_o <= x"d258";
				when 16#01b7# => read_data_o <= x"71e0";
				when 16#01b8# => read_data_o <= x"0050";
				when 16#01b9# => read_data_o <= x"d1e5";
				when 16#01ba# => read_data_o <= x"d1c5";
				when 16#01bb# => read_data_o <= x"d137";
				when 16#01bc# => read_data_o <= x"d1b2";
				when 16#01bd# => read_data_o <= x"d02b";
				when 16#01be# => read_data_o <= x"d0a1";
				when 16#01bf# => read_data_o <= x"d08c";
				when 16#01c0# => read_data_o <= x"d095";
				when 16#01c1# => read_data_o <= x"d095";
				when 16#01c2# => read_data_o <= x"d095";
				when 16#01c3# => read_data_o <= x"d1a8";
				when 16#01c4# => read_data_o <= x"d17f";
				when 16#01c5# => read_data_o <= x"d30c";
				when 16#01c6# => read_data_o <= x"d02b";
				when 16#01c7# => read_data_o <= x"d02b";
				when 16#01c8# => read_data_o <= x"d02b";
				when 16#01c9# => read_data_o <= x"d02b";
				when 16#01ca# => read_data_o <= x"d02b";
				when 16#01cb# => read_data_o <= x"7050";
				when 16#01cc# => read_data_o <= x"0050";
				when 16#01cd# => read_data_o <= x"d14e";
				when 16#01ce# => read_data_o <= x"d160";
				when 16#01cf# => read_data_o <= x"d1b2";
				when 16#01d0# => read_data_o <= x"d1ef";
				when 16#01d1# => read_data_o <= x"d160";
				when 16#01d2# => read_data_o <= x"d1da";
				when 16#01d3# => read_data_o <= x"d02b";
				when 16#01d4# => read_data_o <= x"d0b2";
				when 16#01d5# => read_data_o <= x"d095";
				when 16#01d6# => read_data_o <= x"d095";
				when 16#01d7# => read_data_o <= x"d08c";
				when 16#01d8# => read_data_o <= x"d095";
				when 16#01d9# => read_data_o <= x"d095";
				when 16#01da# => read_data_o <= x"d095";
				when 16#01db# => read_data_o <= x"d1a8";
				when 16#01dc# => read_data_o <= x"d17f";
				when 16#01dd# => read_data_o <= x"d30c";
				when 16#01de# => read_data_o <= x"d02b";
				when 16#01df# => read_data_o <= x"d02b";
				when 16#01e0# => read_data_o <= x"d02b";
				when 16#01e1# => read_data_o <= x"d02b";
				when 16#01e2# => read_data_o <= x"d02b";
				when 16#01e3# => read_data_o <= x"7050";
				when 16#01e4# => read_data_o <= x"02dc";
				when 16#01e5# => read_data_o <= x"d1da";
				when 16#01e6# => read_data_o <= x"d1a2";
				when 16#01e7# => read_data_o <= x"d02b";
				when 16#01e8# => read_data_o <= x"d095";
				when 16#01e9# => read_data_o <= x"d25f";
				when 16#01ea# => read_data_o <= x"d140";
				when 16#01eb# => read_data_o <= x"d2a8";
				when 16#01ec# => read_data_o <= x"d02b";
				when 16#01ed# => read_data_o <= x"d02b";
				when 16#01ee# => read_data_o <= x"d02b";
				when 16#01ef# => read_data_o <= x"d02b";
				when 16#01f0# => read_data_o <= x"d02b";
				when 16#01f1# => read_data_o <= x"d02b";
				when 16#01f2# => read_data_o <= x"7040";
				when 16#01f3# => read_data_o <= x"02fc";
				when 16#01f4# => read_data_o <= x"d02b";
				when 16#01f5# => read_data_o <= x"d137";
				when 16#01f6# => read_data_o <= x"d1ef";
				when 16#01f7# => read_data_o <= x"d1ef";
				when 16#01f8# => read_data_o <= x"d160";
				when 16#01f9# => read_data_o <= x"d1b2";
				when 16#01fa# => read_data_o <= x"d02b";
				when 16#01fb# => read_data_o <= x"d0a1";
				when 16#01fc# => read_data_o <= x"d095";
				when 16#01fd# => read_data_o <= x"d25f";
				when 16#01fe# => read_data_o <= x"d140";
				when 16#01ff# => read_data_o <= x"7110";
				when 16#0200# => read_data_o <= x"02fc";
				when 16#0201# => read_data_o <= x"d02b";
				when 16#0202# => read_data_o <= x"d02b";
				when 16#0203# => read_data_o <= x"d02b";
				when 16#0204# => read_data_o <= x"d02b";
				when 16#0205# => read_data_o <= x"d02b";
				when 16#0206# => read_data_o <= x"d02b";
				when 16#0207# => read_data_o <= x"d02b";
				when 16#0208# => read_data_o <= x"d02b";
				when 16#0209# => read_data_o <= x"7130";
				when 16#020a# => read_data_o <= x"02dc";
				when 16#020b# => read_data_o <= x"d0a1";
				when 16#020c# => read_data_o <= x"d095";
				when 16#020d# => read_data_o <= x"d25f";
				when 16#020e# => read_data_o <= x"d140";
				when 16#020f# => read_data_o <= x"d091";
				when 16#0210# => read_data_o <= x"d02b";
				when 16#0211# => read_data_o <= x"71b0";
				when 16#0212# => read_data_o <= x"02fc";
				when 16#0213# => read_data_o <= x"d1a8";
				when 16#0214# => read_data_o <= x"d198";
				when 16#0215# => read_data_o <= x"d1da";
				when 16#0216# => read_data_o <= x"d02b";
				when 16#0217# => read_data_o <= x"d088";
				when 16#0218# => read_data_o <= x"d0a1";
				when 16#0219# => read_data_o <= x"d095";
				when 16#021a# => read_data_o <= x"d08c";
				when 16#021b# => read_data_o <= x"d0a1";
				when 16#021c# => read_data_o <= x"d0dc";
				when 16#021d# => read_data_o <= x"d25f";
				when 16#021e# => read_data_o <= x"d140";
				when 16#021f# => read_data_o <= x"d2a8";
				when 16#0220# => read_data_o <= x"d02b";
				when 16#0221# => read_data_o <= x"d02b";
				when 16#0222# => read_data_o <= x"d02b";
				when 16#0223# => read_data_o <= x"d02b";
				when 16#0224# => read_data_o <= x"71b0";
				when 16#0225# => read_data_o <= x"02dc";
				when 16#0226# => read_data_o <= x"d0b2";
				when 16#0227# => read_data_o <= x"d095";
				when 16#0228# => read_data_o <= x"d095";
				when 16#0229# => read_data_o <= x"d08c";
				when 16#022a# => read_data_o <= x"d095";
				when 16#022b# => read_data_o <= x"d095";
				when 16#022c# => read_data_o <= x"d0a8";
				when 16#022d# => read_data_o <= x"d1a8";
				when 16#022e# => read_data_o <= x"d17f";
				when 16#022f# => read_data_o <= x"d30c";
				when 16#0230# => read_data_o <= x"d02b";
				when 16#0231# => read_data_o <= x"d02b";
				when 16#0232# => read_data_o <= x"d02b";
				when 16#0233# => read_data_o <= x"d02b";
				when 16#0234# => read_data_o <= x"d02b";
				when 16#0235# => read_data_o <= x"d02b";
				when 16#0236# => read_data_o <= x"d02b";
				when 16#0237# => read_data_o <= x"d02b";
				when 16#0238# => read_data_o <= x"d02b";
				when 16#0239# => read_data_o <= x"7060";
				when 16#023a# => read_data_o <= x"027a";
				when 16#023b# => read_data_o <= x"d02b";
				when 16#023c# => read_data_o <= x"d02b";
				when 16#023d# => read_data_o <= x"d02b";
				when 16#023e# => read_data_o <= x"d02b";
				when 16#023f# => read_data_o <= x"d02b";
				when 16#0240# => read_data_o <= x"d02b";
				when 16#0241# => read_data_o <= x"d02b";
				when 16#0242# => read_data_o <= x"d02b";
				when 16#0243# => read_data_o <= x"d02b";
				when 16#0244# => read_data_o <= x"d02b";
				when 16#0245# => read_data_o <= x"d02b";
				when 16#0246# => read_data_o <= x"d02b";
				when 16#0247# => read_data_o <= x"7040";
				when 16#0248# => read_data_o <= x"022c";
				when 16#0249# => read_data_o <= x"d02b";
				when 16#024a# => read_data_o <= x"7040";
				when 16#024b# => read_data_o <= x"020c";
				when 16#024c# => read_data_o <= x"d02b";
				when 16#024d# => read_data_o <= x"7040";
				when 16#024e# => read_data_o <= x"01ec";
				when 16#024f# => read_data_o <= x"d02b";
				when 16#0250# => read_data_o <= x"7040";
				when 16#0251# => read_data_o <= x"01cc";
				when 16#0252# => read_data_o <= x"d02b";
				when 16#0253# => read_data_o <= x"7040";
				when 16#0254# => read_data_o <= x"01ac";
				when 16#0255# => read_data_o <= x"d02b";
				when 16#0256# => read_data_o <= x"7040";
				when 16#0257# => read_data_o <= x"018c";
				when 16#0258# => read_data_o <= x"d02b";
				when 16#0259# => read_data_o <= x"7040";
				when 16#025a# => read_data_o <= x"016c";
				when 16#025b# => read_data_o <= x"d02b";
				when 16#025c# => read_data_o <= x"7040";
				when 16#025d# => read_data_o <= x"014c";
				when 16#025e# => read_data_o <= x"d02b";
				when 16#025f# => read_data_o <= x"7040";
				when 16#0260# => read_data_o <= x"012c";
				when 16#0261# => read_data_o <= x"d02b";
				when 16#0262# => read_data_o <= x"7040";
				when 16#0263# => read_data_o <= x"010c";
				when 16#0264# => read_data_o <= x"d02b";
				when 16#0265# => read_data_o <= x"ba04";
				when 16#0266# => read_data_o <= x"0000";
				when 16#0267# => read_data_o <= x"0000";
				when 16#0268# => read_data_o <= x"a000";
				when 16#0269# => read_data_o <= x"0270";
				when 16#026a# => read_data_o <= x"d02b";
				when 16#026b# => read_data_o <= x"2404";
				when 16#026c# => read_data_o <= x"7064";
				when 16#026d# => read_data_o <= x"02bc";
				when 16#026e# => read_data_o <= x"a532";
				when 16#026f# => read_data_o <= x"0000";
				when 16#0270# => read_data_o <= x"0000";
				when 16#0271# => read_data_o <= x"0000";
				when 16#0272# => read_data_o <= x"0000";
				when 16#0273# => read_data_o <= x"0000";
				when 16#0274# => read_data_o <= x"0000";
				when 16#0275# => read_data_o <= x"0000";
				when 16#0276# => read_data_o <= x"0000";
				when 16#0277# => read_data_o <= x"0000";
				when 16#0278# => read_data_o <= x"0000";
				when 16#0279# => read_data_o <= x"0000";
				when 16#027a# => read_data_o <= x"0000";
				when 16#027b# => read_data_o <= x"0000";
				when 16#027c# => read_data_o <= x"0000";
				when 16#027d# => read_data_o <= x"0000";
				when 16#027e# => read_data_o <= x"0000";
				when 16#027f# => read_data_o <= x"0000";
				when 16#0280# => read_data_o <= x"0000";
				when 16#0281# => read_data_o <= x"0000";
				when 16#0282# => read_data_o <= x"0000";
				when 16#0283# => read_data_o <= x"0000";
				when 16#0284# => read_data_o <= x"0000";
				when 16#0285# => read_data_o <= x"0000";
				when 16#0286# => read_data_o <= x"0000";
				when 16#0287# => read_data_o <= x"0000";
				when 16#0288# => read_data_o <= x"0000";
				when 16#0289# => read_data_o <= x"0000";
				when 16#028a# => read_data_o <= x"0000";
				when 16#028b# => read_data_o <= x"0000";
				when 16#028c# => read_data_o <= x"0000";
				when 16#028d# => read_data_o <= x"0000";
				when 16#028e# => read_data_o <= x"0000";
				when 16#028f# => read_data_o <= x"0000";
				when 16#0290# => read_data_o <= x"0000";
				when 16#0291# => read_data_o <= x"0000";
				when 16#0292# => read_data_o <= x"0000";
				when 16#0293# => read_data_o <= x"0000";
				when 16#0294# => read_data_o <= x"0000";
				when 16#0295# => read_data_o <= x"0000";
				when 16#0296# => read_data_o <= x"0000";
				when 16#0297# => read_data_o <= x"0000";
				when 16#0298# => read_data_o <= x"0000";
				when 16#0299# => read_data_o <= x"a000";
				when 16#029a# => read_data_o <= x"7064";
				when 16#029b# => read_data_o <= x"02bc";
				when 16#029c# => read_data_o <= x"a58e";
				when 16#029d# => read_data_o <= x"0000";
				when 16#029e# => read_data_o <= x"0000";
				when 16#029f# => read_data_o <= x"0000";
				when 16#02a0# => read_data_o <= x"0000";
				when 16#02a1# => read_data_o <= x"0000";
				when 16#02a2# => read_data_o <= x"0000";
				when 16#02a3# => read_data_o <= x"0000";
				when 16#02a4# => read_data_o <= x"0000";
				when 16#02a5# => read_data_o <= x"0000";
				when 16#02a6# => read_data_o <= x"0000";
				when 16#02a7# => read_data_o <= x"0000";
				when 16#02a8# => read_data_o <= x"0000";
				when 16#02a9# => read_data_o <= x"0000";
				when 16#02aa# => read_data_o <= x"0000";
				when 16#02ab# => read_data_o <= x"0000";
				when 16#02ac# => read_data_o <= x"0000";
				when 16#02ad# => read_data_o <= x"0000";
				when 16#02ae# => read_data_o <= x"0000";
				when 16#02af# => read_data_o <= x"0000";
				when 16#02b0# => read_data_o <= x"0000";
				when 16#02b1# => read_data_o <= x"0000";
				when 16#02b2# => read_data_o <= x"0000";
				when 16#02b3# => read_data_o <= x"0000";
				when 16#02b4# => read_data_o <= x"0000";
				when 16#02b5# => read_data_o <= x"0000";
				when 16#02b6# => read_data_o <= x"0000";
				when 16#02b7# => read_data_o <= x"0000";
				when 16#02b8# => read_data_o <= x"0000";
				when 16#02b9# => read_data_o <= x"0000";
				when 16#02ba# => read_data_o <= x"0000";
				when 16#02bb# => read_data_o <= x"0000";
				when 16#02bc# => read_data_o <= x"0000";
				when 16#02bd# => read_data_o <= x"0000";
				when 16#02be# => read_data_o <= x"0000";
				when 16#02bf# => read_data_o <= x"0000";
				when 16#02c0# => read_data_o <= x"0000";
				when 16#02c1# => read_data_o <= x"0000";
				when 16#02c2# => read_data_o <= x"0000";
				when 16#02c3# => read_data_o <= x"0000";
				when 16#02c4# => read_data_o <= x"0000";
				when 16#02c5# => read_data_o <= x"0000";
				when 16#02c6# => read_data_o <= x"0000";
				when 16#02c7# => read_data_o <= x"a000";
				when 16#02c8# => read_data_o <= x"a592";
				when 16#02c9# => read_data_o <= x"7064";
				when 16#02ca# => read_data_o <= x"0064";
				when 16#02cb# => read_data_o <= x"7064";
				when 16#02cc# => read_data_o <= x"0064";
				when 16#02cd# => read_data_o <= x"5064";
				when 16#02ce# => read_data_o <= x"0190";
				when 16#02cf# => read_data_o <= x"5064";
				when 16#02d0# => read_data_o <= x"02bc";
				when 16#02d1# => read_data_o <= x"70a0";
				when 16#02d2# => read_data_o <= x"02bc";
				when 16#02d3# => read_data_o <= x"50a0";
				when 16#02d4# => read_data_o <= x"0190";
				when 16#02d5# => read_data_o <= x"50a0";
				when 16#02d6# => read_data_o <= x"0064";
				when 16#02d7# => read_data_o <= x"70dc";
				when 16#02d8# => read_data_o <= x"0064";
				when 16#02d9# => read_data_o <= x"50dc";
				when 16#02da# => read_data_o <= x"0190";
				when 16#02db# => read_data_o <= x"50dc";
				when 16#02dc# => read_data_o <= x"02bc";
				when 16#02dd# => read_data_o <= x"7118";
				when 16#02de# => read_data_o <= x"02bc";
				when 16#02df# => read_data_o <= x"5118";
				when 16#02e0# => read_data_o <= x"0190";
				when 16#02e1# => read_data_o <= x"5118";
				when 16#02e2# => read_data_o <= x"0064";
				when 16#02e3# => read_data_o <= x"7154";
				when 16#02e4# => read_data_o <= x"0064";
				when 16#02e5# => read_data_o <= x"5154";
				when 16#02e6# => read_data_o <= x"0190";
				when 16#02e7# => read_data_o <= x"5154";
				when 16#02e8# => read_data_o <= x"02bc";
				when 16#02e9# => read_data_o <= x"7190";
				when 16#02ea# => read_data_o <= x"02bc";
				when 16#02eb# => read_data_o <= x"5190";
				when 16#02ec# => read_data_o <= x"0190";
				when 16#02ed# => read_data_o <= x"5190";
				when 16#02ee# => read_data_o <= x"0064";
				when 16#02ef# => read_data_o <= x"71cc";
				when 16#02f0# => read_data_o <= x"0064";
				when 16#02f1# => read_data_o <= x"51cc";
				when 16#02f2# => read_data_o <= x"0190";
				when 16#02f3# => read_data_o <= x"51cc";
				when 16#02f4# => read_data_o <= x"02bc";
				when 16#02f5# => read_data_o <= x"7208";
				when 16#02f6# => read_data_o <= x"02bc";
				when 16#02f7# => read_data_o <= x"5208";
				when 16#02f8# => read_data_o <= x"0190";
				when 16#02f9# => read_data_o <= x"5208";
				when 16#02fa# => read_data_o <= x"0064";
				when 16#02fb# => read_data_o <= x"7244";
				when 16#02fc# => read_data_o <= x"0064";
				when 16#02fd# => read_data_o <= x"5244";
				when 16#02fe# => read_data_o <= x"0190";
				when 16#02ff# => read_data_o <= x"5244";
				when 16#0300# => read_data_o <= x"02bc";
				when 16#0301# => read_data_o <= x"7280";
				when 16#0302# => read_data_o <= x"02bc";
				when 16#0303# => read_data_o <= x"5280";
				when 16#0304# => read_data_o <= x"0190";
				when 16#0305# => read_data_o <= x"5280";
				when 16#0306# => read_data_o <= x"0064";
				when 16#0307# => read_data_o <= x"72bc";
				when 16#0308# => read_data_o <= x"0064";
				when 16#0309# => read_data_o <= x"52bc";
				when 16#030a# => read_data_o <= x"0190";
				when 16#030b# => read_data_o <= x"52bc";
				when 16#030c# => read_data_o <= x"02bc";
				when 16#030d# => read_data_o <= x"72bc";
				when 16#030e# => read_data_o <= x"02bc";
				when 16#030f# => read_data_o <= x"5190";
				when 16#0310# => read_data_o <= x"02bc";
				when 16#0311# => read_data_o <= x"5064";
				when 16#0312# => read_data_o <= x"02bc";
				when 16#0313# => read_data_o <= x"7064";
				when 16#0314# => read_data_o <= x"0280";
				when 16#0315# => read_data_o <= x"5190";
				when 16#0316# => read_data_o <= x"0280";
				when 16#0317# => read_data_o <= x"52bc";
				when 16#0318# => read_data_o <= x"0280";
				when 16#0319# => read_data_o <= x"72bc";
				when 16#031a# => read_data_o <= x"0244";
				when 16#031b# => read_data_o <= x"5190";
				when 16#031c# => read_data_o <= x"0244";
				when 16#031d# => read_data_o <= x"5064";
				when 16#031e# => read_data_o <= x"0244";
				when 16#031f# => read_data_o <= x"7064";
				when 16#0320# => read_data_o <= x"0208";
				when 16#0321# => read_data_o <= x"5190";
				when 16#0322# => read_data_o <= x"0208";
				when 16#0323# => read_data_o <= x"52bc";
				when 16#0324# => read_data_o <= x"0208";
				when 16#0325# => read_data_o <= x"72bc";
				when 16#0326# => read_data_o <= x"01cc";
				when 16#0327# => read_data_o <= x"5190";
				when 16#0328# => read_data_o <= x"01cc";
				when 16#0329# => read_data_o <= x"5064";
				when 16#032a# => read_data_o <= x"01cc";
				when 16#032b# => read_data_o <= x"7064";
				when 16#032c# => read_data_o <= x"0190";
				when 16#032d# => read_data_o <= x"5190";
				when 16#032e# => read_data_o <= x"0190";
				when 16#032f# => read_data_o <= x"52bc";
				when 16#0330# => read_data_o <= x"0190";
				when 16#0331# => read_data_o <= x"72bc";
				when 16#0332# => read_data_o <= x"0154";
				when 16#0333# => read_data_o <= x"5190";
				when 16#0334# => read_data_o <= x"0154";
				when 16#0335# => read_data_o <= x"5064";
				when 16#0336# => read_data_o <= x"0154";
				when 16#0337# => read_data_o <= x"7064";
				when 16#0338# => read_data_o <= x"0118";
				when 16#0339# => read_data_o <= x"5190";
				when 16#033a# => read_data_o <= x"0118";
				when 16#033b# => read_data_o <= x"52bc";
				when 16#033c# => read_data_o <= x"0118";
				when 16#033d# => read_data_o <= x"72bc";
				when 16#033e# => read_data_o <= x"00dc";
				when 16#033f# => read_data_o <= x"5190";
				when 16#0340# => read_data_o <= x"00dc";
				when 16#0341# => read_data_o <= x"5064";
				when 16#0342# => read_data_o <= x"00dc";
				when 16#0343# => read_data_o <= x"7064";
				when 16#0344# => read_data_o <= x"00a0";
				when 16#0345# => read_data_o <= x"5190";
				when 16#0346# => read_data_o <= x"00a0";
				when 16#0347# => read_data_o <= x"52bc";
				when 16#0348# => read_data_o <= x"00a0";
				when 16#0349# => read_data_o <= x"72bc";
				when 16#034a# => read_data_o <= x"0064";
				when 16#034b# => read_data_o <= x"5190";
				when 16#034c# => read_data_o <= x"0064";
				when 16#034d# => read_data_o <= x"5064";
				when 16#034e# => read_data_o <= x"0064";
				when 16#034f# => read_data_o <= x"a6a0";
				when 16#0350# => read_data_o <= x"2403";
				when 16#0351# => read_data_o <= x"a6e2";
				when 16#0352# => read_data_o <= x"0000";
				when 16#0353# => read_data_o <= x"0000";
				when 16#0354# => read_data_o <= x"0000";
				when 16#0355# => read_data_o <= x"0000";
				when 16#0356# => read_data_o <= x"0000";
				when 16#0357# => read_data_o <= x"0000";
				when 16#0358# => read_data_o <= x"0000";
				when 16#0359# => read_data_o <= x"0000";
				when 16#035a# => read_data_o <= x"0000";
				when 16#035b# => read_data_o <= x"0000";
				when 16#035c# => read_data_o <= x"0000";
				when 16#035d# => read_data_o <= x"0000";
				when 16#035e# => read_data_o <= x"0000";
				when 16#035f# => read_data_o <= x"0000";
				when 16#0360# => read_data_o <= x"0000";
				when 16#0361# => read_data_o <= x"0000";
				when 16#0362# => read_data_o <= x"0000";
				when 16#0363# => read_data_o <= x"0000";
				when 16#0364# => read_data_o <= x"0000";
				when 16#0365# => read_data_o <= x"0000";
				when 16#0366# => read_data_o <= x"0000";
				when 16#0367# => read_data_o <= x"0000";
				when 16#0368# => read_data_o <= x"0000";
				when 16#0369# => read_data_o <= x"0000";
				when 16#036a# => read_data_o <= x"0000";
				when 16#036b# => read_data_o <= x"0000";
				when 16#036c# => read_data_o <= x"0000";
				when 16#036d# => read_data_o <= x"0000";
				when 16#036e# => read_data_o <= x"0000";
				when 16#036f# => read_data_o <= x"0000";
				when 16#0370# => read_data_o <= x"0000";
				when 16#0371# => read_data_o <= x"a000";
				when 16#0372# => read_data_o <= x"027f";
				when 16#0373# => read_data_o <= x"4194";
				when 16#0374# => read_data_o <= x"0285";
				when 16#0375# => read_data_o <= x"4191";
				when 16#0376# => read_data_o <= x"028b";
				when 16#0377# => read_data_o <= x"418e";
				when 16#0378# => read_data_o <= x"0285";
				when 16#0379# => read_data_o <= x"4191";
				when 16#037a# => read_data_o <= x"027f";
				when 16#037b# => read_data_o <= x"4194";
				when 16#037c# => read_data_o <= x"0285";
				when 16#037d# => read_data_o <= x"4191";
				when 16#037e# => read_data_o <= x"028b";
				when 16#037f# => read_data_o <= x"418e";
				when 16#0380# => read_data_o <= x"0285";
				when 16#0381# => read_data_o <= x"4191";
				when 16#0382# => read_data_o <= x"027f";
				when 16#0383# => read_data_o <= x"4194";
				when 16#0384# => read_data_o <= x"0285";
				when 16#0385# => read_data_o <= x"4191";
				when 16#0386# => read_data_o <= x"028b";
				when 16#0387# => read_data_o <= x"418e";
				when 16#0388# => read_data_o <= x"0285";
				when 16#0389# => read_data_o <= x"4191";
				when 16#038a# => read_data_o <= x"027f";
				when 16#038b# => read_data_o <= x"a722";
				when 16#038c# => read_data_o <= x"0000";
				when 16#038d# => read_data_o <= x"0000";
				when 16#038e# => read_data_o <= x"0000";
				when 16#038f# => read_data_o <= x"0000";
				when 16#0390# => read_data_o <= x"0000";
				when 16#0391# => read_data_o <= x"a000";
				when 16#0392# => read_data_o <= x"0000";
				when 16#0393# => read_data_o <= x"0000";
				when 16#0394# => read_data_o <= x"0000";
				when 16#0395# => read_data_o <= x"0000";
				when 16#0396# => read_data_o <= x"0000";
				when 16#0397# => read_data_o <= x"0000";
				when 16#0398# => read_data_o <= x"0000";
				when 16#0399# => read_data_o <= x"0000";
				when 16#039a# => read_data_o <= x"0000";
				when 16#039b# => read_data_o <= x"0000";
				when 16#039c# => read_data_o <= x"0000";
				when 16#039d# => read_data_o <= x"0000";
				when 16#039e# => read_data_o <= x"0000";
				when 16#039f# => read_data_o <= x"0000";
				when 16#03a0# => read_data_o <= x"0000";
				when 16#03a1# => read_data_o <= x"0000";
				when 16#03a2# => read_data_o <= x"0000";
				when 16#03a3# => read_data_o <= x"0000";
				when 16#03a4# => read_data_o <= x"0000";
				when 16#03a5# => read_data_o <= x"0000";
				when 16#03a6# => read_data_o <= x"0000";
				when 16#03a7# => read_data_o <= x"0000";
				when 16#03a8# => read_data_o <= x"0000";
				when 16#03a9# => read_data_o <= x"0000";
				when 16#03aa# => read_data_o <= x"0000";
				when 16#03ab# => read_data_o <= x"0000";
				when 16#03ac# => read_data_o <= x"0000";
				when 16#03ad# => read_data_o <= x"0000";
				when 16#03ae# => read_data_o <= x"0000";
				when 16#03af# => read_data_o <= x"0000";
				when 16#03b0# => read_data_o <= x"0000";
				when 16#03b1# => read_data_o <= x"a000";
				when 16#03b2# => read_data_o <= x"0000";
				when 16#03b3# => read_data_o <= x"0000";
				when 16#03b4# => read_data_o <= x"0000";
				when 16#03b5# => read_data_o <= x"0000";
				when 16#03b6# => read_data_o <= x"0000";
				when 16#03b7# => read_data_o <= x"0000";
				when 16#03b8# => read_data_o <= x"0000";
				when 16#03b9# => read_data_o <= x"0000";
				when 16#03ba# => read_data_o <= x"0000";
				when 16#03bb# => read_data_o <= x"0000";
				when 16#03bc# => read_data_o <= x"0000";
				when 16#03bd# => read_data_o <= x"0000";
				when 16#03be# => read_data_o <= x"0000";
				when 16#03bf# => read_data_o <= x"0000";
				when 16#03c0# => read_data_o <= x"0000";
				when 16#03c1# => read_data_o <= x"0000";
				when 16#03c2# => read_data_o <= x"0000";
				when 16#03c3# => read_data_o <= x"0000";
				when 16#03c4# => read_data_o <= x"0000";
				when 16#03c5# => read_data_o <= x"0000";
				when 16#03c6# => read_data_o <= x"0000";
				when 16#03c7# => read_data_o <= x"0000";
				when 16#03c8# => read_data_o <= x"0000";
				when 16#03c9# => read_data_o <= x"0000";
				when 16#03ca# => read_data_o <= x"0000";
				when 16#03cb# => read_data_o <= x"0000";
				when 16#03cc# => read_data_o <= x"0000";
				when 16#03cd# => read_data_o <= x"0000";
				when 16#03ce# => read_data_o <= x"0000";
				when 16#03cf# => read_data_o <= x"0000";
				when 16#03d0# => read_data_o <= x"0000";
				when 16#03d1# => read_data_o <= x"a000";
				when 16#03d2# => read_data_o <= x"0000";
				when 16#03d3# => read_data_o <= x"0000";
				when 16#03d4# => read_data_o <= x"0000";
				when 16#03d5# => read_data_o <= x"0000";
				when 16#03d6# => read_data_o <= x"0000";
				when 16#03d7# => read_data_o <= x"0000";
				when 16#03d8# => read_data_o <= x"0000";
				when 16#03d9# => read_data_o <= x"0000";
				when 16#03da# => read_data_o <= x"0000";
				when 16#03db# => read_data_o <= x"0000";
				when 16#03dc# => read_data_o <= x"0000";
				when 16#03dd# => read_data_o <= x"0000";
				when 16#03de# => read_data_o <= x"0000";
				when 16#03df# => read_data_o <= x"0000";
				when 16#03e0# => read_data_o <= x"0000";
				when 16#03e1# => read_data_o <= x"0000";
				when 16#03e2# => read_data_o <= x"0000";
				when 16#03e3# => read_data_o <= x"0000";
				when 16#03e4# => read_data_o <= x"0000";
				when 16#03e5# => read_data_o <= x"0000";
				when 16#03e6# => read_data_o <= x"0000";
				when 16#03e7# => read_data_o <= x"0000";
				when 16#03e8# => read_data_o <= x"0000";
				when 16#03e9# => read_data_o <= x"0000";
				when 16#03ea# => read_data_o <= x"0000";
				when 16#03eb# => read_data_o <= x"0000";
				when 16#03ec# => read_data_o <= x"0000";
				when 16#03ed# => read_data_o <= x"0000";
				when 16#03ee# => read_data_o <= x"0000";
				when 16#03ef# => read_data_o <= x"0000";
				when 16#03f0# => read_data_o <= x"0000";
				when 16#03f1# => read_data_o <= x"a000";
				when 16#03f2# => read_data_o <= x"7064";
				when 16#03f3# => read_data_o <= x"00ba";
				when 16#03f4# => read_data_o <= x"0064";
				when 16#03f5# => read_data_o <= x"00b7";
				when 16#03f6# => read_data_o <= x"0064";
				when 16#03f7# => read_data_o <= x"00b5";
				when 16#03f8# => read_data_o <= x"006c";
				when 16#03f9# => read_data_o <= x"00b7";
				when 16#03fa# => read_data_o <= x"006b";
				when 16#03fb# => read_data_o <= x"00bb";
				when 16#03fc# => read_data_o <= x"0064";
				when 16#03fd# => read_data_o <= x"00b5";
				when 16#03fe# => read_data_o <= x"0064";
				when 16#03ff# => read_data_o <= x"00b7";
				when 16#0400# => read_data_o <= x"0064";
				when 16#0401# => read_data_o <= x"00b7";
				when 16#0402# => read_data_o <= x"0064";
				when 16#0403# => read_data_o <= x"00b7";
				when 16#0404# => read_data_o <= x"0064";
				when 16#0405# => read_data_o <= x"00c0";
				when 16#0406# => read_data_o <= x"0064";
				when 16#0407# => read_data_o <= x"00b7";
				when 16#0408# => read_data_o <= x"0064";
				when 16#0409# => read_data_o <= x"00b6";
				when 16#040a# => read_data_o <= x"0064";
				when 16#040b# => read_data_o <= x"00b9";
				when 16#040c# => read_data_o <= x"0064";
				when 16#040d# => read_data_o <= x"00ba";
				when 16#040e# => read_data_o <= x"0064";
				when 16#040f# => read_data_o <= x"00bc";
				when 16#0410# => read_data_o <= x"0064";
				when 16#0411# => read_data_o <= x"00bc";
				when 16#0412# => read_data_o <= x"0064";
				when 16#0413# => read_data_o <= x"00b8";
				when 16#0414# => read_data_o <= x"006b";
				when 16#0415# => read_data_o <= x"00b9";
				when 16#0416# => read_data_o <= x"0069";
				when 16#0417# => read_data_o <= x"00b4";
				when 16#0418# => read_data_o <= x"0064";
				when 16#0419# => read_data_o <= x"00b0";
				when 16#041a# => read_data_o <= x"0064";
				when 16#041b# => read_data_o <= x"00b3";
				when 16#041c# => read_data_o <= x"006b";
				when 16#041d# => read_data_o <= x"00b6";
				when 16#041e# => read_data_o <= x"0064";
				when 16#041f# => read_data_o <= x"00bd";
				when 16#0420# => read_data_o <= x"0064";
				when 16#0421# => read_data_o <= x"00b6";
				when 16#0422# => read_data_o <= x"0064";
				when 16#0423# => read_data_o <= x"00b8";
				when 16#0424# => read_data_o <= x"006b";
				when 16#0425# => read_data_o <= x"00ba";
				when 16#0426# => read_data_o <= x"0064";
				when 16#0427# => read_data_o <= x"00ba";
				when 16#0428# => read_data_o <= x"0064";
				when 16#0429# => read_data_o <= x"00b5";
				when 16#042a# => read_data_o <= x"0064";
				when 16#042b# => read_data_o <= x"00b9";
				when 16#042c# => read_data_o <= x"0064";
				when 16#042d# => read_data_o <= x"00b1";
				when 16#042e# => read_data_o <= x"0064";
				when 16#042f# => read_data_o <= x"00c2";
				when 16#0430# => read_data_o <= x"0064";
				when 16#0431# => read_data_o <= x"00b9";
				when 16#0432# => read_data_o <= x"0064";
				when 16#0433# => read_data_o <= x"00b9";
				when 16#0434# => read_data_o <= x"0064";
				when 16#0435# => read_data_o <= x"00b9";
				when 16#0436# => read_data_o <= x"0064";
				when 16#0437# => read_data_o <= x"00bd";
				when 16#0438# => read_data_o <= x"0064";
				when 16#0439# => read_data_o <= x"00bb";
				when 16#043a# => read_data_o <= x"0064";
				when 16#043b# => read_data_o <= x"00bf";
				when 16#043c# => read_data_o <= x"0065";
				when 16#043d# => read_data_o <= x"00b8";
				when 16#043e# => read_data_o <= x"0064";
				when 16#043f# => read_data_o <= x"00bf";
				when 16#0440# => read_data_o <= x"0064";
				when 16#0441# => read_data_o <= x"00b8";
				when 16#0442# => read_data_o <= x"0064";
				when 16#0443# => read_data_o <= x"00be";
				when 16#0444# => read_data_o <= x"0064";
				when 16#0445# => read_data_o <= x"00b4";
				when 16#0446# => read_data_o <= x"0064";
				when 16#0447# => read_data_o <= x"00bb";
				when 16#0448# => read_data_o <= x"0072";
				when 16#0449# => read_data_o <= x"00b6";
				when 16#044a# => read_data_o <= x"0064";
				when 16#044b# => read_data_o <= x"00bd";
				when 16#044c# => read_data_o <= x"0064";
				when 16#044d# => read_data_o <= x"00bc";
				when 16#044e# => read_data_o <= x"0064";
				when 16#044f# => read_data_o <= x"00b8";
				when 16#0450# => read_data_o <= x"006a";
				when 16#0451# => read_data_o <= x"00b6";
				when 16#0452# => read_data_o <= x"0064";
				when 16#0453# => read_data_o <= x"00bc";
				when 16#0454# => read_data_o <= x"0064";
				when 16#0455# => read_data_o <= x"00be";
				when 16#0456# => read_data_o <= x"0064";
				when 16#0457# => read_data_o <= x"00be";
				when 16#0458# => read_data_o <= x"0064";
				when 16#0459# => read_data_o <= x"00b5";
				when 16#045a# => read_data_o <= x"0064";
				when 16#045b# => read_data_o <= x"00bd";
				when 16#045c# => read_data_o <= x"0065";
				when 16#045d# => read_data_o <= x"00ba";
				when 16#045e# => read_data_o <= x"0064";
				when 16#045f# => read_data_o <= x"00b8";
				when 16#0460# => read_data_o <= x"0064";
				when 16#0461# => read_data_o <= x"00c2";
				when 16#0462# => read_data_o <= x"0064";
				when 16#0463# => read_data_o <= x"00c6";
				when 16#0464# => read_data_o <= x"0064";
				when 16#0465# => read_data_o <= x"00d1";
				when 16#0466# => read_data_o <= x"0081";
				when 16#0467# => read_data_o <= x"00cb";
				when 16#0468# => read_data_o <= x"0072";
				when 16#0469# => read_data_o <= x"00ca";
				when 16#046a# => read_data_o <= x"006d";
				when 16#046b# => read_data_o <= x"00bd";
				when 16#046c# => read_data_o <= x"0066";
				when 16#046d# => read_data_o <= x"00b7";
				when 16#046e# => read_data_o <= x"0064";
				when 16#046f# => read_data_o <= x"00b5";
				when 16#0470# => read_data_o <= x"0064";
				when 16#0471# => read_data_o <= x"00ba";
				when 16#0472# => read_data_o <= x"0064";
				when 16#0473# => read_data_o <= x"00b3";
				when 16#0474# => read_data_o <= x"0064";
				when 16#0475# => read_data_o <= x"00b2";
				when 16#0476# => read_data_o <= x"0064";
				when 16#0477# => read_data_o <= x"00b6";
				when 16#0478# => read_data_o <= x"0068";
				when 16#0479# => read_data_o <= x"00c1";
				when 16#047a# => read_data_o <= x"0064";
				when 16#047b# => read_data_o <= x"00b5";
				when 16#047c# => read_data_o <= x"006c";
				when 16#047d# => read_data_o <= x"00b7";
				when 16#047e# => read_data_o <= x"0064";
				when 16#047f# => read_data_o <= x"00be";
				when 16#0480# => read_data_o <= x"0064";
				when 16#0481# => read_data_o <= x"00bb";
				when 16#0482# => read_data_o <= x"0064";
				when 16#0483# => read_data_o <= x"00c1";
				when 16#0484# => read_data_o <= x"0066";
				when 16#0485# => read_data_o <= x"00b8";
				when 16#0486# => read_data_o <= x"0064";
				when 16#0487# => read_data_o <= x"00b7";
				when 16#0488# => read_data_o <= x"0069";
				when 16#0489# => read_data_o <= x"00b9";
				when 16#048a# => read_data_o <= x"0067";
				when 16#048b# => read_data_o <= x"00c1";
				when 16#048c# => read_data_o <= x"0064";
				when 16#048d# => read_data_o <= x"00bc";
				when 16#048e# => read_data_o <= x"0064";
				when 16#048f# => read_data_o <= x"00c0";
				when 16#0490# => read_data_o <= x"0064";
				when 16#0491# => read_data_o <= x"00bc";
				when 16#0492# => read_data_o <= x"0064";
				when 16#0493# => read_data_o <= x"00c2";
				when 16#0494# => read_data_o <= x"0068";
				when 16#0495# => read_data_o <= x"00bd";
				when 16#0496# => read_data_o <= x"0069";
				when 16#0497# => read_data_o <= x"00c1";
				when 16#0498# => read_data_o <= x"0064";
				when 16#0499# => read_data_o <= x"00bf";
				when 16#049a# => read_data_o <= x"006d";
				when 16#049b# => read_data_o <= x"00b9";
				when 16#049c# => read_data_o <= x"0064";
				when 16#049d# => read_data_o <= x"00bb";
				when 16#049e# => read_data_o <= x"0064";
				when 16#049f# => read_data_o <= x"00cb";
				when 16#04a0# => read_data_o <= x"0064";
				when 16#04a1# => read_data_o <= x"00b8";
				when 16#04a2# => read_data_o <= x"0064";
				when 16#04a3# => read_data_o <= x"00b6";
				when 16#04a4# => read_data_o <= x"0064";
				when 16#04a5# => read_data_o <= x"00be";
				when 16#04a6# => read_data_o <= x"0064";
				when 16#04a7# => read_data_o <= x"00b8";
				when 16#04a8# => read_data_o <= x"006f";
				when 16#04a9# => read_data_o <= x"00ba";
				when 16#04aa# => read_data_o <= x"0064";
				when 16#04ab# => read_data_o <= x"00b7";
				when 16#04ac# => read_data_o <= x"0067";
				when 16#04ad# => read_data_o <= x"00ba";
				when 16#04ae# => read_data_o <= x"0067";
				when 16#04af# => read_data_o <= x"00c4";
				when 16#04b0# => read_data_o <= x"0064";
				when 16#04b1# => read_data_o <= x"00bb";
				when 16#04b2# => read_data_o <= x"0064";
				when 16#04b3# => read_data_o <= x"00be";
				when 16#04b4# => read_data_o <= x"0064";
				when 16#04b5# => read_data_o <= x"00b7";
				when 16#04b6# => read_data_o <= x"0064";
				when 16#04b7# => read_data_o <= x"00ba";
				when 16#04b8# => read_data_o <= x"0064";
				when 16#04b9# => read_data_o <= x"00be";
				when 16#04ba# => read_data_o <= x"0068";
				when 16#04bb# => read_data_o <= x"00bc";
				when 16#04bc# => read_data_o <= x"0064";
				when 16#04bd# => read_data_o <= x"00bd";
				when 16#04be# => read_data_o <= x"0064";
				when 16#04bf# => read_data_o <= x"00be";
				when 16#04c0# => read_data_o <= x"0064";
				when 16#04c1# => read_data_o <= x"00bf";
				when 16#04c2# => read_data_o <= x"0064";
				when 16#04c3# => read_data_o <= x"00bb";
				when 16#04c4# => read_data_o <= x"0064";
				when 16#04c5# => read_data_o <= x"00bb";
				when 16#04c6# => read_data_o <= x"0066";
				when 16#04c7# => read_data_o <= x"00ba";
				when 16#04c8# => read_data_o <= x"0064";
				when 16#04c9# => read_data_o <= x"00bc";
				when 16#04ca# => read_data_o <= x"0068";
				when 16#04cb# => read_data_o <= x"00bf";
				when 16#04cc# => read_data_o <= x"006e";
				when 16#04cd# => read_data_o <= x"00c4";
				when 16#04ce# => read_data_o <= x"006c";
				when 16#04cf# => read_data_o <= x"00c0";
				when 16#04d0# => read_data_o <= x"0064";
				when 16#04d1# => read_data_o <= x"00bf";
				when 16#04d2# => read_data_o <= x"0064";
				when 16#04d3# => read_data_o <= x"00c5";
				when 16#04d4# => read_data_o <= x"0064";
				when 16#04d5# => read_data_o <= x"00c7";
				when 16#04d6# => read_data_o <= x"0070";
				when 16#04d7# => read_data_o <= x"00bb";
				when 16#04d8# => read_data_o <= x"0064";
				when 16#04d9# => read_data_o <= x"00c6";
				when 16#04da# => read_data_o <= x"0065";
				when 16#04db# => read_data_o <= x"00be";
				when 16#04dc# => read_data_o <= x"0065";
				when 16#04dd# => read_data_o <= x"00cb";
				when 16#04de# => read_data_o <= x"0064";
				when 16#04df# => read_data_o <= x"00bf";
				when 16#04e0# => read_data_o <= x"0064";
				when 16#04e1# => read_data_o <= x"00c1";
				when 16#04e2# => read_data_o <= x"2069";
				when 16#04e3# => read_data_o <= x"20bf";
				when 16#04e4# => read_data_o <= x"2064";
				when 16#04e5# => read_data_o <= x"20ca";
				when 16#04e6# => read_data_o <= x"2069";
				when 16#04e7# => read_data_o <= x"00cb";
				when 16#04e8# => read_data_o <= x"006b";
				when 16#04e9# => read_data_o <= x"00c3";
				when 16#04ea# => read_data_o <= x"0064";
				when 16#04eb# => read_data_o <= x"00c7";
				when 16#04ec# => read_data_o <= x"0064";
				when 16#04ed# => read_data_o <= x"00c2";
				when 16#04ee# => read_data_o <= x"0064";
				when 16#04ef# => read_data_o <= x"00c5";
				when 16#04f0# => read_data_o <= x"0076";
				when 16#04f1# => read_data_o <= x"00c9";
				when 16#04f2# => read_data_o <= x"006b";
				when 16#04f3# => read_data_o <= x"00cd";
				when 16#04f4# => read_data_o <= x"007a";
				when 16#04f5# => read_data_o <= x"00c6";
				when 16#04f6# => read_data_o <= x"0087";
				when 16#04f7# => read_data_o <= x"00d5";
				when 16#04f8# => read_data_o <= x"00a5";
				when 16#04f9# => read_data_o <= x"00d7";
				when 16#04fa# => read_data_o <= x"00b6";
				when 16#04fb# => read_data_o <= x"00dc";
				when 16#04fc# => read_data_o <= x"00ca";
				when 16#04fd# => read_data_o <= x"00ea";
				when 16#04fe# => read_data_o <= x"00dc";
				when 16#04ff# => read_data_o <= x"00fc";
				when 16#0500# => read_data_o <= x"0102";
				when 16#0501# => read_data_o <= x"010d";
				when 16#0502# => read_data_o <= x"0116";
				when 16#0503# => read_data_o <= x"0120";
				when 16#0504# => read_data_o <= x"012a";
				when 16#0505# => read_data_o <= x"0134";
				when 16#0506# => read_data_o <= x"013f";
				when 16#0507# => read_data_o <= x"014a";
				when 16#0508# => read_data_o <= x"0155";
				when 16#0509# => read_data_o <= x"0161";
				when 16#050a# => read_data_o <= x"016d";
				when 16#050b# => read_data_o <= x"0179";
				when 16#050c# => read_data_o <= x"0185";
				when 16#050d# => read_data_o <= x"0192";
				when 16#050e# => read_data_o <= x"019f";
				when 16#050f# => read_data_o <= x"01ac";
				when 16#0510# => read_data_o <= x"01ba";
				when 16#0511# => read_data_o <= x"01c8";
				when 16#0512# => read_data_o <= x"01d6";
				when 16#0513# => read_data_o <= x"01e4";
				when 16#0514# => read_data_o <= x"01f3";
				when 16#0515# => read_data_o <= x"0202";
				when 16#0516# => read_data_o <= x"0211";
				when 16#0517# => read_data_o <= x"0220";
				when 16#0518# => read_data_o <= x"0230";
				when 16#0519# => read_data_o <= x"023f";
				when 16#051a# => read_data_o <= x"024e";
				when 16#051b# => read_data_o <= x"025c";
				when 16#051c# => read_data_o <= x"0269";
				when 16#051d# => read_data_o <= x"0273";
				when 16#051e# => read_data_o <= x"027b";
				when 16#051f# => read_data_o <= x"027e";
				when 16#0520# => read_data_o <= x"027f";
				when 16#0521# => read_data_o <= x"027d";
				when 16#0522# => read_data_o <= x"0278";
				when 16#0523# => read_data_o <= x"026f";
				when 16#0524# => read_data_o <= x"0263";
				when 16#0525# => read_data_o <= x"0256";
				when 16#0526# => read_data_o <= x"0247";
				when 16#0527# => read_data_o <= x"0238";
				when 16#0528# => read_data_o <= x"0229";
				when 16#0529# => read_data_o <= x"0219";
				when 16#052a# => read_data_o <= x"020a";
				when 16#052b# => read_data_o <= x"01fb";
				when 16#052c# => read_data_o <= x"01ec";
				when 16#052d# => read_data_o <= x"01dd";
				when 16#052e# => read_data_o <= x"01cf";
				when 16#052f# => read_data_o <= x"01c0";
				when 16#0530# => read_data_o <= x"01b3";
				when 16#0531# => read_data_o <= x"01a5";
				when 16#0532# => read_data_o <= x"0198";
				when 16#0533# => read_data_o <= x"018b";
				when 16#0534# => read_data_o <= x"017e";
				when 16#0535# => read_data_o <= x"0172";
				when 16#0536# => read_data_o <= x"0166";
				when 16#0537# => read_data_o <= x"015a";
				when 16#0538# => read_data_o <= x"014f";
				when 16#0539# => read_data_o <= x"0144";
				when 16#053a# => read_data_o <= x"0139";
				when 16#053b# => read_data_o <= x"012f";
				when 16#053c# => read_data_o <= x"0125";
				when 16#053d# => read_data_o <= x"011b";
				when 16#053e# => read_data_o <= x"0110";
				when 16#053f# => read_data_o <= x"0108";
				when 16#0540# => read_data_o <= x"00ee";
				when 16#0541# => read_data_o <= x"00ff";
				when 16#0542# => read_data_o <= x"00db";
				when 16#0543# => read_data_o <= x"00f0";
				when 16#0544# => read_data_o <= x"00c7";
				when 16#0545# => read_data_o <= x"00df";
				when 16#0546# => read_data_o <= x"00b3";
				when 16#0547# => read_data_o <= x"00d9";
				when 16#0548# => read_data_o <= x"00a1";
				when 16#0549# => read_data_o <= x"00d3";
				when 16#054a# => read_data_o <= x"0094";
				when 16#054b# => read_data_o <= x"00d2";
				when 16#054c# => read_data_o <= x"0082";
				when 16#054d# => read_data_o <= x"00cc";
				when 16#054e# => read_data_o <= x"006c";
				when 16#054f# => read_data_o <= x"00ca";
				when 16#0550# => read_data_o <= x"0069";
				when 16#0551# => read_data_o <= x"00cd";
				when 16#0552# => read_data_o <= x"006d";
				when 16#0553# => read_data_o <= x"00ca";
				when 16#0554# => read_data_o <= x"006a";
				when 16#0555# => read_data_o <= x"00cf";
				when 16#0556# => read_data_o <= x"0068";
				when 16#0557# => read_data_o <= x"00bb";
				when 16#0558# => read_data_o <= x"0064";
				when 16#0559# => read_data_o <= x"00c6";
				when 16#055a# => read_data_o <= x"0069";
				when 16#055b# => read_data_o <= x"00c5";
				when 16#055c# => read_data_o <= x"0072";
				when 16#055d# => read_data_o <= x"00c8";
				when 16#055e# => read_data_o <= x"0064";
				when 16#055f# => read_data_o <= x"00c5";
				when 16#0560# => read_data_o <= x"0064";
				when 16#0561# => read_data_o <= x"00cb";
				when 16#0562# => read_data_o <= x"0064";
				when 16#0563# => read_data_o <= x"00c2";
				when 16#0564# => read_data_o <= x"0064";
				when 16#0565# => read_data_o <= x"00bf";
				when 16#0566# => read_data_o <= x"0064";
				when 16#0567# => read_data_o <= x"00bf";
				when 16#0568# => read_data_o <= x"0075";
				when 16#0569# => read_data_o <= x"00bd";
				when 16#056a# => read_data_o <= x"0064";
				when 16#056b# => read_data_o <= x"00c4";
				when 16#056c# => read_data_o <= x"0064";
				when 16#056d# => read_data_o <= x"00c5";
				when 16#056e# => read_data_o <= x"0064";
				when 16#056f# => read_data_o <= x"00c8";
				when 16#0570# => read_data_o <= x"0064";
				when 16#0571# => read_data_o <= x"00bd";
				when 16#0572# => read_data_o <= x"0064";
				when 16#0573# => read_data_o <= x"00c7";
				when 16#0574# => read_data_o <= x"0064";
				when 16#0575# => read_data_o <= x"00c3";
				when 16#0576# => read_data_o <= x"0064";
				when 16#0577# => read_data_o <= x"00c3";
				when 16#0578# => read_data_o <= x"0067";
				when 16#0579# => read_data_o <= x"00bd";
				when 16#057a# => read_data_o <= x"0064";
				when 16#057b# => read_data_o <= x"00c5";
				when 16#057c# => read_data_o <= x"0064";
				when 16#057d# => read_data_o <= x"00c3";
				when 16#057e# => read_data_o <= x"0064";
				when 16#057f# => read_data_o <= x"00ba";
				when 16#0580# => read_data_o <= x"006d";
				when 16#0581# => read_data_o <= x"00b7";
				when 16#0582# => read_data_o <= x"0064";
				when 16#0583# => read_data_o <= x"00bf";
				when 16#0584# => read_data_o <= x"0067";
				when 16#0585# => read_data_o <= x"00bb";
				when 16#0586# => read_data_o <= x"0064";
				when 16#0587# => read_data_o <= x"00bc";
				when 16#0588# => read_data_o <= x"0064";
				when 16#0589# => read_data_o <= x"00ba";
				when 16#058a# => read_data_o <= x"0071";
				when 16#058b# => read_data_o <= x"00be";
				when 16#058c# => read_data_o <= x"0064";
				when 16#058d# => read_data_o <= x"00bd";
				when 16#058e# => read_data_o <= x"0072";
				when 16#058f# => read_data_o <= x"00bc";
				when 16#0590# => read_data_o <= x"0064";
				when 16#0591# => read_data_o <= x"00b5";
				when 16#0592# => read_data_o <= x"0064";
				when 16#0593# => read_data_o <= x"00bd";
				when 16#0594# => read_data_o <= x"0064";
				when 16#0595# => read_data_o <= x"00bc";
				when 16#0596# => read_data_o <= x"0064";
				when 16#0597# => read_data_o <= x"00b5";
				when 16#0598# => read_data_o <= x"0069";
				when 16#0599# => read_data_o <= x"00b7";
				when 16#059a# => read_data_o <= x"0064";
				when 16#059b# => read_data_o <= x"00bb";
				when 16#059c# => read_data_o <= x"0064";
				when 16#059d# => read_data_o <= x"00bd";
				when 16#059e# => read_data_o <= x"0068";
				when 16#059f# => read_data_o <= x"00b5";
				when 16#05a0# => read_data_o <= x"0064";
				when 16#05a1# => read_data_o <= x"00c1";
				when 16#05a2# => read_data_o <= x"0064";
				when 16#05a3# => read_data_o <= x"00b7";
				when 16#05a4# => read_data_o <= x"0064";
				when 16#05a5# => read_data_o <= x"00b4";
				when 16#05a6# => read_data_o <= x"0064";
				when 16#05a7# => read_data_o <= x"00bd";
				when 16#05a8# => read_data_o <= x"0064";
				when 16#05a9# => read_data_o <= x"00b4";
				when 16#05aa# => read_data_o <= x"0064";
				when 16#05ab# => read_data_o <= x"00c0";
				when 16#05ac# => read_data_o <= x"0064";
				when 16#05ad# => read_data_o <= x"00cc";
				when 16#05ae# => read_data_o <= x"0064";
				when 16#05af# => read_data_o <= x"00c4";
				when 16#05b0# => read_data_o <= x"0064";
				when 16#05b1# => read_data_o <= x"00c2";
				when 16#05b2# => read_data_o <= x"0068";
				when 16#05b3# => read_data_o <= x"00b7";
				when 16#05b4# => read_data_o <= x"0064";
				when 16#05b5# => read_data_o <= x"00ba";
				when 16#05b6# => read_data_o <= x"0064";
				when 16#05b7# => read_data_o <= x"00b8";
				when 16#05b8# => read_data_o <= x"0064";
				when 16#05b9# => read_data_o <= x"00ba";
				when 16#05ba# => read_data_o <= x"006b";
				when 16#05bb# => read_data_o <= x"00b2";
				when 16#05bc# => read_data_o <= x"0064";
				when 16#05bd# => read_data_o <= x"00bf";
				when 16#05be# => read_data_o <= x"0067";
				when 16#05bf# => read_data_o <= x"00b7";
				when 16#05c0# => read_data_o <= x"0066";
				when 16#05c1# => read_data_o <= x"00bb";
				when 16#05c2# => read_data_o <= x"006a";
				when 16#05c3# => read_data_o <= x"00b4";
				when 16#05c4# => read_data_o <= x"0064";
				when 16#05c5# => read_data_o <= x"00bc";
				when 16#05c6# => read_data_o <= x"0064";
				when 16#05c7# => read_data_o <= x"00bd";
				when 16#05c8# => read_data_o <= x"0064";
				when 16#05c9# => read_data_o <= x"00b7";
				when 16#05ca# => read_data_o <= x"0064";
				when 16#05cb# => read_data_o <= x"00bc";
				when 16#05cc# => read_data_o <= x"0064";
				when 16#05cd# => read_data_o <= x"00bb";
				when 16#05ce# => read_data_o <= x"0064";
				when 16#05cf# => read_data_o <= x"00bc";
				when 16#05d0# => read_data_o <= x"0064";
				when 16#05d1# => read_data_o <= x"00b9";
				when 16#05d2# => read_data_o <= x"0064";
				when 16#05d3# => read_data_o <= x"00bd";
				when 16#05d4# => read_data_o <= x"0067";
				when 16#05d5# => read_data_o <= x"00c3";
				when 16#05d6# => read_data_o <= x"0067";
				when 16#05d7# => read_data_o <= x"00ce";
				when 16#05d8# => read_data_o <= x"0066";
				when 16#05d9# => read_data_o <= x"00d8";
				when 16#05da# => read_data_o <= x"007c";
				when 16#05db# => read_data_o <= x"00d1";
				when 16#05dc# => read_data_o <= x"006e";
				when 16#05dd# => read_data_o <= x"00c5";
				when 16#05de# => read_data_o <= x"0064";
				when 16#05df# => read_data_o <= x"00c6";
				when 16#05e0# => read_data_o <= x"0064";
				when 16#05e1# => read_data_o <= x"00bc";
				when 16#05e2# => read_data_o <= x"0064";
				when 16#05e3# => read_data_o <= x"00b8";
				when 16#05e4# => read_data_o <= x"0064";
				when 16#05e5# => read_data_o <= x"00ba";
				when 16#05e6# => read_data_o <= x"0064";
				when 16#05e7# => read_data_o <= x"00b7";
				when 16#05e8# => read_data_o <= x"0069";
				when 16#05e9# => read_data_o <= x"00bb";
				when 16#05ea# => read_data_o <= x"0064";
				when 16#05eb# => read_data_o <= x"00b9";
				when 16#05ec# => read_data_o <= x"0064";
				when 16#05ed# => read_data_o <= x"00c0";
				when 16#05ee# => read_data_o <= x"0068";
				when 16#05ef# => read_data_o <= x"00bc";
				when 16#05f0# => read_data_o <= x"0064";
				when 16#05f1# => read_data_o <= x"00be";
				when 16#05f2# => read_data_o <= x"0064";
				when 16#05f3# => read_data_o <= x"00b3";
				when 16#05f4# => read_data_o <= x"0064";
				when 16#05f5# => read_data_o <= x"00bd";
				when 16#05f6# => read_data_o <= x"0064";
				when 16#05f7# => read_data_o <= x"00b7";
				when 16#05f8# => read_data_o <= x"0067";
				when 16#05f9# => read_data_o <= x"00be";
				when 16#05fa# => read_data_o <= x"0064";
				when 16#05fb# => read_data_o <= x"00b8";
				when 16#05fc# => read_data_o <= x"0064";
				when 16#05fd# => read_data_o <= x"00b8";
				when 16#05fe# => read_data_o <= x"0064";
				when 16#05ff# => read_data_o <= x"00b3";
				when 16#0600# => read_data_o <= x"0064";
				when 16#0601# => read_data_o <= x"00b7";
				when 16#0602# => read_data_o <= x"0064";
				when 16#0603# => read_data_o <= x"00b8";
				when 16#0604# => read_data_o <= x"0064";
				when 16#0605# => read_data_o <= x"00b8";
				when 16#0606# => read_data_o <= x"0064";
				when 16#0607# => read_data_o <= x"00c5";
				when 16#0608# => read_data_o <= x"0064";
				when 16#0609# => read_data_o <= x"00c4";
				when 16#060a# => read_data_o <= x"0064";
				when 16#060b# => read_data_o <= x"00ba";
				when 16#060c# => read_data_o <= x"006f";
				when 16#060d# => read_data_o <= x"00c1";
				when 16#060e# => read_data_o <= x"0066";
				when 16#060f# => read_data_o <= x"00bf";
				when 16#0610# => read_data_o <= x"0069";
				when 16#0611# => read_data_o <= x"00b8";
				when 16#0612# => read_data_o <= x"0069";
				when 16#0613# => read_data_o <= x"00b7";
				when 16#0614# => read_data_o <= x"0069";
				when 16#0615# => read_data_o <= x"00b8";
				when 16#0616# => read_data_o <= x"0064";
				when 16#0617# => read_data_o <= x"00b2";
				when 16#0618# => read_data_o <= x"0064";
				when 16#0619# => read_data_o <= x"00b9";
				when 16#061a# => read_data_o <= x"0064";
				when 16#061b# => read_data_o <= x"00bc";
				when 16#061c# => read_data_o <= x"0064";
				when 16#061d# => read_data_o <= x"00b4";
				when 16#061e# => read_data_o <= x"0067";
				when 16#061f# => read_data_o <= x"00b6";
				when 16#0620# => read_data_o <= x"0064";
				when 16#0621# => read_data_o <= x"00c1";
				when 16#0622# => read_data_o <= x"0064";
				when 16#0623# => read_data_o <= x"00bb";
				when 16#0624# => read_data_o <= x"0064";
				when 16#0625# => read_data_o <= x"00b5";
				when 16#0626# => read_data_o <= x"0069";
				when 16#0627# => read_data_o <= x"00b3";
				when 16#0628# => read_data_o <= x"0064";
				when 16#0629# => read_data_o <= x"00b4";
				when 16#062a# => read_data_o <= x"0064";
				when 16#062b# => read_data_o <= x"00bb";
				when 16#062c# => read_data_o <= x"0064";
				when 16#062d# => read_data_o <= x"00ba";
				when 16#062e# => read_data_o <= x"0065";
				when 16#062f# => read_data_o <= x"00c5";
				when 16#0630# => read_data_o <= x"0064";
				when 16#0631# => read_data_o <= x"00b8";
				when 16#0632# => read_data_o <= x"0064";
				when 16#0633# => read_data_o <= x"00ba";
				when 16#0634# => read_data_o <= x"006a";
				when 16#0635# => read_data_o <= x"00ba";
				when 16#0636# => read_data_o <= x"0064";
				when 16#0637# => read_data_o <= x"00bc";
				when 16#0638# => read_data_o <= x"0064";
				when 16#0639# => read_data_o <= x"00b9";
				when 16#063a# => read_data_o <= x"0064";
				when 16#063b# => read_data_o <= x"00b5";
				when 16#063c# => read_data_o <= x"0064";
				when 16#063d# => read_data_o <= x"00b6";
				when 16#063e# => read_data_o <= x"0064";
				when 16#063f# => read_data_o <= x"00b4";
				when 16#0640# => read_data_o <= x"0064";
				when 16#0641# => read_data_o <= x"00bb";
				when 16#0642# => read_data_o <= x"0064";
				when 16#0643# => read_data_o <= x"00bf";
				when 16#0644# => read_data_o <= x"006b";
				when 16#0645# => read_data_o <= x"00bc";
				when 16#0646# => read_data_o <= x"0064";
				when 16#0647# => read_data_o <= x"00bf";
				when 16#0648# => read_data_o <= x"0064";
				when 16#0649# => read_data_o <= x"00b9";
				when 16#064a# => read_data_o <= x"0064";
				when 16#064b# => read_data_o <= x"00b7";
				when 16#064c# => read_data_o <= x"2000";
				when 16#064d# => read_data_o <= x"2000";
				when 16#064e# => read_data_o <= x"2000";
				when 16#064f# => read_data_o <= x"2000";
				when 16#0650# => read_data_o <= x"2000";
				when 16#0651# => read_data_o <= x"2405";
				when 16#0652# => read_data_o <= x"7064";
				when 16#0653# => read_data_o <= x"3064";
				when 16#0654# => read_data_o <= x"3064";
				when 16#0655# => read_data_o <= x"3064";
				when 16#0656# => read_data_o <= x"3064";
				when 16#0657# => read_data_o <= x"3064";
				when 16#0658# => read_data_o <= x"3064";
				when 16#0659# => read_data_o <= x"3064";
				when 16#065a# => read_data_o <= x"3064";
				when 16#065b# => read_data_o <= x"3064";
				when 16#065c# => read_data_o <= x"3064";
				when 16#065d# => read_data_o <= x"3064";
				when 16#065e# => read_data_o <= x"3064";
				when 16#065f# => read_data_o <= x"3064";
				when 16#0660# => read_data_o <= x"3064";
				when 16#0661# => read_data_o <= x"3064";
				when 16#0662# => read_data_o <= x"3064";
				when 16#0663# => read_data_o <= x"3064";
				when 16#0664# => read_data_o <= x"3064";
				when 16#0665# => read_data_o <= x"3064";
				when 16#0666# => read_data_o <= x"3064";
				when 16#0667# => read_data_o <= x"3064";
				when 16#0668# => read_data_o <= x"3064";
				when 16#0669# => read_data_o <= x"3064";
				when 16#066a# => read_data_o <= x"3064";
				when 16#066b# => read_data_o <= x"3064";
				when 16#066c# => read_data_o <= x"3064";
				when 16#066d# => read_data_o <= x"3064";
				when 16#066e# => read_data_o <= x"3064";
				when 16#066f# => read_data_o <= x"3064";
				when 16#0670# => read_data_o <= x"3064";
				when 16#0671# => read_data_o <= x"3064";
				when 16#0672# => read_data_o <= x"3064";
				when 16#0673# => read_data_o <= x"3064";
				when 16#0674# => read_data_o <= x"3064";
				when 16#0675# => read_data_o <= x"3064";
				when 16#0676# => read_data_o <= x"3064";
				when 16#0677# => read_data_o <= x"3064";
				when 16#0678# => read_data_o <= x"3064";
				when 16#0679# => read_data_o <= x"3064";
				when 16#067a# => read_data_o <= x"3064";
				when 16#067b# => read_data_o <= x"3064";
				when 16#067c# => read_data_o <= x"3064";
				when 16#067d# => read_data_o <= x"3064";
				when 16#067e# => read_data_o <= x"3064";
				when 16#067f# => read_data_o <= x"3064";
				when 16#0680# => read_data_o <= x"3064";
				when 16#0681# => read_data_o <= x"3064";
				when 16#0682# => read_data_o <= x"3064";
				when 16#0683# => read_data_o <= x"3064";
				when 16#0684# => read_data_o <= x"3064";
				when 16#0685# => read_data_o <= x"3064";
				when 16#0686# => read_data_o <= x"3064";
				when 16#0687# => read_data_o <= x"3064";
				when 16#0688# => read_data_o <= x"3064";
				when 16#0689# => read_data_o <= x"3064";
				when 16#068a# => read_data_o <= x"3064";
				when 16#068b# => read_data_o <= x"3064";
				when 16#068c# => read_data_o <= x"3064";
				when 16#068d# => read_data_o <= x"3064";
				when 16#068e# => read_data_o <= x"3064";
				when 16#068f# => read_data_o <= x"3064";
				when 16#0690# => read_data_o <= x"3064";
				when 16#0691# => read_data_o <= x"3064";
				when 16#0692# => read_data_o <= x"3064";
				when 16#0693# => read_data_o <= x"3064";
				when 16#0694# => read_data_o <= x"3064";
				when 16#0695# => read_data_o <= x"3064";
				when 16#0696# => read_data_o <= x"3064";
				when 16#0697# => read_data_o <= x"3064";
				when 16#0698# => read_data_o <= x"3064";
				when 16#0699# => read_data_o <= x"3064";
				when 16#069a# => read_data_o <= x"3064";
				when 16#069b# => read_data_o <= x"3064";
				when 16#069c# => read_data_o <= x"3064";
				when 16#069d# => read_data_o <= x"3064";
				when 16#069e# => read_data_o <= x"3064";
				when 16#069f# => read_data_o <= x"3064";
				when 16#06a0# => read_data_o <= x"3064";
				when 16#06a1# => read_data_o <= x"3064";
				when 16#06a2# => read_data_o <= x"3064";
				when 16#06a3# => read_data_o <= x"3064";
				when 16#06a4# => read_data_o <= x"3064";
				when 16#06a5# => read_data_o <= x"3064";
				when 16#06a6# => read_data_o <= x"3064";
				when 16#06a7# => read_data_o <= x"3064";
				when 16#06a8# => read_data_o <= x"3064";
				when 16#06a9# => read_data_o <= x"3064";
				when 16#06aa# => read_data_o <= x"3064";
				when 16#06ab# => read_data_o <= x"3064";
				when 16#06ac# => read_data_o <= x"3064";
				when 16#06ad# => read_data_o <= x"3064";
				when 16#06ae# => read_data_o <= x"3064";
				when 16#06af# => read_data_o <= x"3064";
				when 16#06b0# => read_data_o <= x"3064";
				when 16#06b1# => read_data_o <= x"3064";
				when 16#06b2# => read_data_o <= x"3064";
				when 16#06b3# => read_data_o <= x"3064";
				when 16#06b4# => read_data_o <= x"3064";
				when 16#06b5# => read_data_o <= x"3064";
				when 16#06b6# => read_data_o <= x"3064";
				when 16#06b7# => read_data_o <= x"3064";
				when 16#06b8# => read_data_o <= x"3064";
				when 16#06b9# => read_data_o <= x"3064";
				when 16#06ba# => read_data_o <= x"3064";
				when 16#06bb# => read_data_o <= x"3064";
				when 16#06bc# => read_data_o <= x"3064";
				when 16#06bd# => read_data_o <= x"3064";
				when 16#06be# => read_data_o <= x"3064";
				when 16#06bf# => read_data_o <= x"3064";
				when 16#06c0# => read_data_o <= x"3064";
				when 16#06c1# => read_data_o <= x"3064";
				when 16#06c2# => read_data_o <= x"3064";
				when 16#06c3# => read_data_o <= x"3064";
				when 16#06c4# => read_data_o <= x"3064";
				when 16#06c5# => read_data_o <= x"3064";
				when 16#06c6# => read_data_o <= x"3064";
				when 16#06c7# => read_data_o <= x"3064";
				when 16#06c8# => read_data_o <= x"3064";
				when 16#06c9# => read_data_o <= x"3064";
				when 16#06ca# => read_data_o <= x"3064";
				when 16#06cb# => read_data_o <= x"3064";
				when 16#06cc# => read_data_o <= x"3064";
				when 16#06cd# => read_data_o <= x"3064";
				when 16#06ce# => read_data_o <= x"3064";
				when 16#06cf# => read_data_o <= x"3064";
				when 16#06d0# => read_data_o <= x"3064";
				when 16#06d1# => read_data_o <= x"3064";
				when 16#06d2# => read_data_o <= x"3064";
				when 16#06d3# => read_data_o <= x"3064";
				when 16#06d4# => read_data_o <= x"3064";
				when 16#06d5# => read_data_o <= x"3064";
				when 16#06d6# => read_data_o <= x"3064";
				when 16#06d7# => read_data_o <= x"3064";
				when 16#06d8# => read_data_o <= x"3064";
				when 16#06d9# => read_data_o <= x"3064";
				when 16#06da# => read_data_o <= x"3064";
				when 16#06db# => read_data_o <= x"3064";
				when 16#06dc# => read_data_o <= x"3064";
				when 16#06dd# => read_data_o <= x"3064";
				when 16#06de# => read_data_o <= x"3064";
				when 16#06df# => read_data_o <= x"3064";
				when 16#06e0# => read_data_o <= x"3064";
				when 16#06e1# => read_data_o <= x"3064";
				when 16#06e2# => read_data_o <= x"3064";
				when 16#06e3# => read_data_o <= x"3064";
				when 16#06e4# => read_data_o <= x"3064";
				when 16#06e5# => read_data_o <= x"3064";
				when 16#06e6# => read_data_o <= x"3064";
				when 16#06e7# => read_data_o <= x"3064";
				when 16#06e8# => read_data_o <= x"3064";
				when 16#06e9# => read_data_o <= x"3064";
				when 16#06ea# => read_data_o <= x"3064";
				when 16#06eb# => read_data_o <= x"3064";
				when 16#06ec# => read_data_o <= x"3064";
				when 16#06ed# => read_data_o <= x"3064";
				when 16#06ee# => read_data_o <= x"3064";
				when 16#06ef# => read_data_o <= x"3064";
				when 16#06f0# => read_data_o <= x"3064";
				when 16#06f1# => read_data_o <= x"3064";
				when 16#06f2# => read_data_o <= x"3064";
				when 16#06f3# => read_data_o <= x"3064";
				when 16#06f4# => read_data_o <= x"3064";
				when 16#06f5# => read_data_o <= x"3064";
				when 16#06f6# => read_data_o <= x"3064";
				when 16#06f7# => read_data_o <= x"3064";
				when 16#06f8# => read_data_o <= x"3064";
				when 16#06f9# => read_data_o <= x"3064";
				when 16#06fa# => read_data_o <= x"3064";
				when 16#06fb# => read_data_o <= x"3064";
				when 16#06fc# => read_data_o <= x"3064";
				when 16#06fd# => read_data_o <= x"3064";
				when 16#06fe# => read_data_o <= x"3064";
				when 16#06ff# => read_data_o <= x"3064";
				when 16#0700# => read_data_o <= x"3064";
				when 16#0701# => read_data_o <= x"3064";
				when 16#0702# => read_data_o <= x"3064";
				when 16#0703# => read_data_o <= x"3064";
				when 16#0704# => read_data_o <= x"3064";
				when 16#0705# => read_data_o <= x"3064";
				when 16#0706# => read_data_o <= x"3064";
				when 16#0707# => read_data_o <= x"3064";
				when 16#0708# => read_data_o <= x"3064";
				when 16#0709# => read_data_o <= x"3064";
				when 16#070a# => read_data_o <= x"3064";
				when 16#070b# => read_data_o <= x"3064";
				when 16#070c# => read_data_o <= x"3064";
				when 16#070d# => read_data_o <= x"3064";
				when 16#070e# => read_data_o <= x"3064";
				when 16#070f# => read_data_o <= x"3064";
				when 16#0710# => read_data_o <= x"3064";
				when 16#0711# => read_data_o <= x"3064";
				when 16#0712# => read_data_o <= x"3064";
				when 16#0713# => read_data_o <= x"3064";
				when 16#0714# => read_data_o <= x"3064";
				when 16#0715# => read_data_o <= x"3064";
				when 16#0716# => read_data_o <= x"3064";
				when 16#0717# => read_data_o <= x"3064";
				when 16#0718# => read_data_o <= x"3064";
				when 16#0719# => read_data_o <= x"3064";
				when 16#071a# => read_data_o <= x"3064";
				when 16#071b# => read_data_o <= x"3064";
				when 16#071c# => read_data_o <= x"3064";
				when 16#071d# => read_data_o <= x"3064";
				when 16#071e# => read_data_o <= x"3064";
				when 16#071f# => read_data_o <= x"3064";
				when 16#0720# => read_data_o <= x"3064";
				when 16#0721# => read_data_o <= x"3064";
				when 16#0722# => read_data_o <= x"3064";
				when 16#0723# => read_data_o <= x"3064";
				when 16#0724# => read_data_o <= x"3064";
				when 16#0725# => read_data_o <= x"3064";
				when 16#0726# => read_data_o <= x"3064";
				when 16#0727# => read_data_o <= x"3064";
				when 16#0728# => read_data_o <= x"3064";
				when 16#0729# => read_data_o <= x"3064";
				when 16#072a# => read_data_o <= x"3064";
				when 16#072b# => read_data_o <= x"3064";
				when 16#072c# => read_data_o <= x"3064";
				when 16#072d# => read_data_o <= x"3064";
				when 16#072e# => read_data_o <= x"3064";
				when 16#072f# => read_data_o <= x"3064";
				when 16#0730# => read_data_o <= x"3064";
				when 16#0731# => read_data_o <= x"3064";
				when 16#0732# => read_data_o <= x"3064";
				when 16#0733# => read_data_o <= x"3064";
				when 16#0734# => read_data_o <= x"3064";
				when 16#0735# => read_data_o <= x"3064";
				when 16#0736# => read_data_o <= x"3064";
				when 16#0737# => read_data_o <= x"3064";
				when 16#0738# => read_data_o <= x"3064";
				when 16#0739# => read_data_o <= x"3064";
				when 16#073a# => read_data_o <= x"3064";
				when 16#073b# => read_data_o <= x"3064";
				when 16#073c# => read_data_o <= x"3064";
				when 16#073d# => read_data_o <= x"3064";
				when 16#073e# => read_data_o <= x"3064";
				when 16#073f# => read_data_o <= x"3064";
				when 16#0740# => read_data_o <= x"3064";
				when 16#0741# => read_data_o <= x"3064";
				when 16#0742# => read_data_o <= x"3064";
				when 16#0743# => read_data_o <= x"3064";
				when 16#0744# => read_data_o <= x"3064";
				when 16#0745# => read_data_o <= x"3064";
				when 16#0746# => read_data_o <= x"3064";
				when 16#0747# => read_data_o <= x"3064";
				when 16#0748# => read_data_o <= x"3064";
				when 16#0749# => read_data_o <= x"3064";
				when 16#074a# => read_data_o <= x"3064";
				when 16#074b# => read_data_o <= x"3064";
				when 16#074c# => read_data_o <= x"3064";
				when 16#074d# => read_data_o <= x"3064";
				when 16#074e# => read_data_o <= x"3064";
				when 16#074f# => read_data_o <= x"3064";
				when 16#0750# => read_data_o <= x"3064";
				when 16#0751# => read_data_o <= x"3064";
				when 16#0752# => read_data_o <= x"3064";
				when 16#0753# => read_data_o <= x"3064";
				when 16#0754# => read_data_o <= x"3064";
				when 16#0755# => read_data_o <= x"3064";
				when 16#0756# => read_data_o <= x"3064";
				when 16#0757# => read_data_o <= x"3064";
				when 16#0758# => read_data_o <= x"3064";
				when 16#0759# => read_data_o <= x"3064";
				when 16#075a# => read_data_o <= x"3064";
				when 16#075b# => read_data_o <= x"3064";
				when 16#075c# => read_data_o <= x"3064";
				when 16#075d# => read_data_o <= x"3064";
				when 16#075e# => read_data_o <= x"3064";
				when 16#075f# => read_data_o <= x"3064";
				when 16#0760# => read_data_o <= x"3064";
				when 16#0761# => read_data_o <= x"3064";
				when 16#0762# => read_data_o <= x"3064";
				when 16#0763# => read_data_o <= x"3064";
				when 16#0764# => read_data_o <= x"3064";
				when 16#0765# => read_data_o <= x"3064";
				when 16#0766# => read_data_o <= x"3064";
				when 16#0767# => read_data_o <= x"3064";
				when 16#0768# => read_data_o <= x"3064";
				when 16#0769# => read_data_o <= x"3064";
				when 16#076a# => read_data_o <= x"3064";
				when 16#076b# => read_data_o <= x"3064";
				when 16#076c# => read_data_o <= x"3064";
				when 16#076d# => read_data_o <= x"3064";
				when 16#076e# => read_data_o <= x"3064";
				when 16#076f# => read_data_o <= x"3064";
				when 16#0770# => read_data_o <= x"3064";
				when 16#0771# => read_data_o <= x"3064";
				when 16#0772# => read_data_o <= x"3064";
				when 16#0773# => read_data_o <= x"3064";
				when 16#0774# => read_data_o <= x"3064";
				when 16#0775# => read_data_o <= x"3064";
				when 16#0776# => read_data_o <= x"3064";
				when 16#0777# => read_data_o <= x"3064";
				when 16#0778# => read_data_o <= x"3064";
				when 16#0779# => read_data_o <= x"3064";
				when 16#077a# => read_data_o <= x"3064";
				when 16#077b# => read_data_o <= x"3064";
				when 16#077c# => read_data_o <= x"3064";
				when 16#077d# => read_data_o <= x"3064";
				when 16#077e# => read_data_o <= x"3064";
				when 16#077f# => read_data_o <= x"3064";
				when 16#0780# => read_data_o <= x"3064";
				when 16#0781# => read_data_o <= x"3064";
				when 16#0782# => read_data_o <= x"3064";
				when 16#0783# => read_data_o <= x"3064";
				when 16#0784# => read_data_o <= x"3064";
				when 16#0785# => read_data_o <= x"3064";
				when 16#0786# => read_data_o <= x"3064";
				when 16#0787# => read_data_o <= x"3064";
				when 16#0788# => read_data_o <= x"3064";
				when 16#0789# => read_data_o <= x"3064";
				when 16#078a# => read_data_o <= x"3064";
				when 16#078b# => read_data_o <= x"3064";
				when 16#078c# => read_data_o <= x"3064";
				when 16#078d# => read_data_o <= x"3064";
				when 16#078e# => read_data_o <= x"3064";
				when 16#078f# => read_data_o <= x"3064";
				when 16#0790# => read_data_o <= x"3064";
				when 16#0791# => read_data_o <= x"3064";
				when 16#0792# => read_data_o <= x"3064";
				when 16#0793# => read_data_o <= x"3064";
				when 16#0794# => read_data_o <= x"3064";
				when 16#0795# => read_data_o <= x"3064";
				when 16#0796# => read_data_o <= x"3064";
				when 16#0797# => read_data_o <= x"3064";
				when 16#0798# => read_data_o <= x"3064";
				when 16#0799# => read_data_o <= x"3064";
				when 16#079a# => read_data_o <= x"3064";
				when 16#079b# => read_data_o <= x"3064";
				when 16#079c# => read_data_o <= x"3064";
				when 16#079d# => read_data_o <= x"3064";
				when 16#079e# => read_data_o <= x"3064";
				when 16#079f# => read_data_o <= x"3064";
				when 16#07a0# => read_data_o <= x"3064";
				when 16#07a1# => read_data_o <= x"3064";
				when 16#07a2# => read_data_o <= x"3064";
				when 16#07a3# => read_data_o <= x"3064";
				when 16#07a4# => read_data_o <= x"3064";
				when 16#07a5# => read_data_o <= x"3064";
				when 16#07a6# => read_data_o <= x"3064";
				when 16#07a7# => read_data_o <= x"3064";
				when 16#07a8# => read_data_o <= x"3064";
				when 16#07a9# => read_data_o <= x"3064";
				when 16#07aa# => read_data_o <= x"3064";
				when 16#07ab# => read_data_o <= x"3064";
				when 16#07ac# => read_data_o <= x"3064";
				when 16#07ad# => read_data_o <= x"3064";
				when 16#07ae# => read_data_o <= x"3064";
				when 16#07af# => read_data_o <= x"3064";
				when 16#07b0# => read_data_o <= x"3064";
				when 16#07b1# => read_data_o <= x"3064";
				when 16#07b2# => read_data_o <= x"3064";
				when 16#07b3# => read_data_o <= x"3064";
				when 16#07b4# => read_data_o <= x"3064";
				when 16#07b5# => read_data_o <= x"3064";
				when 16#07b6# => read_data_o <= x"3064";
				when 16#07b7# => read_data_o <= x"3064";
				when 16#07b8# => read_data_o <= x"3064";
				when 16#07b9# => read_data_o <= x"3064";
				when 16#07ba# => read_data_o <= x"3064";
				when 16#07bb# => read_data_o <= x"3064";
				when 16#07bc# => read_data_o <= x"3064";
				when 16#07bd# => read_data_o <= x"3064";
				when 16#07be# => read_data_o <= x"3064";
				when 16#07bf# => read_data_o <= x"3064";
				when 16#07c0# => read_data_o <= x"3064";
				when 16#07c1# => read_data_o <= x"3064";
				when 16#07c2# => read_data_o <= x"3064";
				when 16#07c3# => read_data_o <= x"3064";
				when 16#07c4# => read_data_o <= x"3064";
				when 16#07c5# => read_data_o <= x"3064";
				when 16#07c6# => read_data_o <= x"3064";
				when 16#07c7# => read_data_o <= x"3064";
				when 16#07c8# => read_data_o <= x"3064";
				when 16#07c9# => read_data_o <= x"3064";
				when 16#07ca# => read_data_o <= x"3064";
				when 16#07cb# => read_data_o <= x"3064";
				when 16#07cc# => read_data_o <= x"3064";
				when 16#07cd# => read_data_o <= x"3064";
				when 16#07ce# => read_data_o <= x"3064";
				when 16#07cf# => read_data_o <= x"3064";
				when 16#07d0# => read_data_o <= x"3064";
				when 16#07d1# => read_data_o <= x"3064";
				when 16#07d2# => read_data_o <= x"3064";
				when 16#07d3# => read_data_o <= x"3064";
				when 16#07d4# => read_data_o <= x"3064";
				when 16#07d5# => read_data_o <= x"3064";
				when 16#07d6# => read_data_o <= x"3064";
				when 16#07d7# => read_data_o <= x"3064";
				when 16#07d8# => read_data_o <= x"3064";
				when 16#07d9# => read_data_o <= x"3064";
				when 16#07da# => read_data_o <= x"3064";
				when 16#07db# => read_data_o <= x"3064";
				when 16#07dc# => read_data_o <= x"3064";
				when 16#07dd# => read_data_o <= x"3064";
				when 16#07de# => read_data_o <= x"3064";
				when 16#07df# => read_data_o <= x"3064";
				when 16#07e0# => read_data_o <= x"3064";
				when 16#07e1# => read_data_o <= x"3064";
				when 16#07e2# => read_data_o <= x"3064";
				when 16#07e3# => read_data_o <= x"3064";
				when 16#07e4# => read_data_o <= x"3064";
				when 16#07e5# => read_data_o <= x"3064";
				when 16#07e6# => read_data_o <= x"3064";
				when 16#07e7# => read_data_o <= x"3064";
				when 16#07e8# => read_data_o <= x"3064";
				when 16#07e9# => read_data_o <= x"3064";
				when 16#07ea# => read_data_o <= x"3064";
				when 16#07eb# => read_data_o <= x"3064";
				when 16#07ec# => read_data_o <= x"3064";
				when 16#07ed# => read_data_o <= x"3064";
				when 16#07ee# => read_data_o <= x"3064";
				when 16#07ef# => read_data_o <= x"3064";
				when 16#07f0# => read_data_o <= x"3064";
				when 16#07f1# => read_data_o <= x"3064";
				when 16#07f2# => read_data_o <= x"3064";
				when 16#07f3# => read_data_o <= x"3064";
				when 16#07f4# => read_data_o <= x"3064";
				when 16#07f5# => read_data_o <= x"3064";
				when 16#07f6# => read_data_o <= x"3064";
				when 16#07f7# => read_data_o <= x"3064";
				when 16#07f8# => read_data_o <= x"3064";
				when 16#07f9# => read_data_o <= x"3064";
				when 16#07fa# => read_data_o <= x"3064";
				when 16#07fb# => read_data_o <= x"3064";
				when 16#07fc# => read_data_o <= x"3064";
				when 16#07fd# => read_data_o <= x"3064";
				when 16#07fe# => read_data_o <= x"3064";
				when 16#07ff# => read_data_o <= x"3064";
				when 16#0800# => read_data_o <= x"3064";
				when 16#0801# => read_data_o <= x"3064";
				when 16#0802# => read_data_o <= x"3064";
				when 16#0803# => read_data_o <= x"3064";
				when 16#0804# => read_data_o <= x"3064";
				when 16#0805# => read_data_o <= x"3064";
				when 16#0806# => read_data_o <= x"3064";
				when 16#0807# => read_data_o <= x"3064";
				when 16#0808# => read_data_o <= x"3064";
				when 16#0809# => read_data_o <= x"3064";
				when 16#080a# => read_data_o <= x"3064";
				when 16#080b# => read_data_o <= x"3064";
				when 16#080c# => read_data_o <= x"3064";
				when 16#080d# => read_data_o <= x"3064";
				when 16#080e# => read_data_o <= x"3064";
				when 16#080f# => read_data_o <= x"3064";
				when 16#0810# => read_data_o <= x"3064";
				when 16#0811# => read_data_o <= x"3064";
				when 16#0812# => read_data_o <= x"3064";
				when 16#0813# => read_data_o <= x"3064";
				when 16#0814# => read_data_o <= x"3064";
				when 16#0815# => read_data_o <= x"3064";
				when 16#0816# => read_data_o <= x"3064";
				when 16#0817# => read_data_o <= x"3064";
				when 16#0818# => read_data_o <= x"3064";
				when 16#0819# => read_data_o <= x"3064";
				when 16#081a# => read_data_o <= x"3064";
				when 16#081b# => read_data_o <= x"3064";
				when 16#081c# => read_data_o <= x"3064";
				when 16#081d# => read_data_o <= x"3064";
				when 16#081e# => read_data_o <= x"3064";
				when 16#081f# => read_data_o <= x"3064";
				when 16#0820# => read_data_o <= x"3064";
				when 16#0821# => read_data_o <= x"3064";
				when 16#0822# => read_data_o <= x"3064";
				when 16#0823# => read_data_o <= x"3064";
				when 16#0824# => read_data_o <= x"3064";
				when 16#0825# => read_data_o <= x"3064";
				when 16#0826# => read_data_o <= x"3064";
				when 16#0827# => read_data_o <= x"3064";
				when 16#0828# => read_data_o <= x"3064";
				when 16#0829# => read_data_o <= x"3064";
				when 16#082a# => read_data_o <= x"3064";
				when 16#082b# => read_data_o <= x"3064";
				when 16#082c# => read_data_o <= x"3064";
				when 16#082d# => read_data_o <= x"3064";
				when 16#082e# => read_data_o <= x"3064";
				when 16#082f# => read_data_o <= x"3064";
				when 16#0830# => read_data_o <= x"3064";
				when 16#0831# => read_data_o <= x"3064";
				when 16#0832# => read_data_o <= x"3064";
				when 16#0833# => read_data_o <= x"3064";
				when 16#0834# => read_data_o <= x"3064";
				when 16#0835# => read_data_o <= x"3064";
				when 16#0836# => read_data_o <= x"3064";
				when 16#0837# => read_data_o <= x"3064";
				when 16#0838# => read_data_o <= x"3064";
				when 16#0839# => read_data_o <= x"3064";
				when 16#083a# => read_data_o <= x"3064";
				when 16#083b# => read_data_o <= x"3064";
				when 16#083c# => read_data_o <= x"3064";
				when 16#083d# => read_data_o <= x"3064";
				when 16#083e# => read_data_o <= x"3064";
				when 16#083f# => read_data_o <= x"3064";
				when 16#0840# => read_data_o <= x"3064";
				when 16#0841# => read_data_o <= x"3064";
				when 16#0842# => read_data_o <= x"3064";
				when 16#0843# => read_data_o <= x"3064";
				when 16#0844# => read_data_o <= x"3064";
				when 16#0845# => read_data_o <= x"3064";
				when 16#0846# => read_data_o <= x"3064";
				when 16#0847# => read_data_o <= x"3064";
				when 16#0848# => read_data_o <= x"3064";
				when 16#0849# => read_data_o <= x"3064";
				when 16#084a# => read_data_o <= x"3064";
				when 16#084b# => read_data_o <= x"3064";
				when 16#084c# => read_data_o <= x"3064";
				when 16#084d# => read_data_o <= x"3064";
				when 16#084e# => read_data_o <= x"3064";
				when 16#084f# => read_data_o <= x"3064";
				when 16#0850# => read_data_o <= x"3064";
				when 16#0851# => read_data_o <= x"3064";
				when 16#0852# => read_data_o <= x"3064";
				when 16#0853# => read_data_o <= x"3064";
				when 16#0854# => read_data_o <= x"3064";
				when 16#0855# => read_data_o <= x"3064";
				when 16#0856# => read_data_o <= x"3064";
				when 16#0857# => read_data_o <= x"3064";
				when 16#0858# => read_data_o <= x"3064";
				when 16#0859# => read_data_o <= x"3064";
				when 16#085a# => read_data_o <= x"3064";
				when 16#085b# => read_data_o <= x"3064";
				when 16#085c# => read_data_o <= x"3064";
				when 16#085d# => read_data_o <= x"3064";
				when 16#085e# => read_data_o <= x"3064";
				when 16#085f# => read_data_o <= x"3064";
				when 16#0860# => read_data_o <= x"3064";
				when 16#0861# => read_data_o <= x"3064";
				when 16#0862# => read_data_o <= x"3064";
				when 16#0863# => read_data_o <= x"3064";
				when 16#0864# => read_data_o <= x"3064";
				when 16#0865# => read_data_o <= x"3064";
				when 16#0866# => read_data_o <= x"3064";
				when 16#0867# => read_data_o <= x"3064";
				when 16#0868# => read_data_o <= x"3064";
				when 16#0869# => read_data_o <= x"3064";
				when 16#086a# => read_data_o <= x"3064";
				when 16#086b# => read_data_o <= x"3064";
				when 16#086c# => read_data_o <= x"3064";
				when 16#086d# => read_data_o <= x"3064";
				when 16#086e# => read_data_o <= x"3064";
				when 16#086f# => read_data_o <= x"3064";
				when 16#0870# => read_data_o <= x"3064";
				when 16#0871# => read_data_o <= x"3064";
				when 16#0872# => read_data_o <= x"3064";
				when 16#0873# => read_data_o <= x"3064";
				when 16#0874# => read_data_o <= x"3064";
				when 16#0875# => read_data_o <= x"3064";
				when 16#0876# => read_data_o <= x"3064";
				when 16#0877# => read_data_o <= x"3064";
				when 16#0878# => read_data_o <= x"3064";
				when 16#0879# => read_data_o <= x"3064";
				when 16#087a# => read_data_o <= x"3064";
				when 16#087b# => read_data_o <= x"3064";
				when 16#087c# => read_data_o <= x"3064";
				when 16#087d# => read_data_o <= x"3064";
				when 16#087e# => read_data_o <= x"3064";
				when 16#087f# => read_data_o <= x"3064";
				when 16#0880# => read_data_o <= x"3064";
				when 16#0881# => read_data_o <= x"3064";
				when 16#0882# => read_data_o <= x"3064";
				when 16#0883# => read_data_o <= x"3064";
				when 16#0884# => read_data_o <= x"3064";
				when 16#0885# => read_data_o <= x"3064";
				when 16#0886# => read_data_o <= x"3064";
				when 16#0887# => read_data_o <= x"3064";
				when 16#0888# => read_data_o <= x"3064";
				when 16#0889# => read_data_o <= x"3064";
				when 16#088a# => read_data_o <= x"3064";
				when 16#088b# => read_data_o <= x"3064";
				when 16#088c# => read_data_o <= x"3064";
				when 16#088d# => read_data_o <= x"3064";
				when 16#088e# => read_data_o <= x"3064";
				when 16#088f# => read_data_o <= x"3064";
				when 16#0890# => read_data_o <= x"3064";
				when 16#0891# => read_data_o <= x"3064";
				when 16#0892# => read_data_o <= x"3064";
				when 16#0893# => read_data_o <= x"3064";
				when 16#0894# => read_data_o <= x"3064";
				when 16#0895# => read_data_o <= x"3064";
				when 16#0896# => read_data_o <= x"3064";
				when 16#0897# => read_data_o <= x"3064";
				when 16#0898# => read_data_o <= x"3064";
				when 16#0899# => read_data_o <= x"3064";
				when 16#089a# => read_data_o <= x"3064";
				when 16#089b# => read_data_o <= x"3064";
				when 16#089c# => read_data_o <= x"3064";
				when 16#089d# => read_data_o <= x"3064";
				when 16#089e# => read_data_o <= x"3064";
				when 16#089f# => read_data_o <= x"3064";
				when 16#08a0# => read_data_o <= x"3064";
				when 16#08a1# => read_data_o <= x"3064";
				when 16#08a2# => read_data_o <= x"3064";
				when 16#08a3# => read_data_o <= x"3064";
				when 16#08a4# => read_data_o <= x"3064";
				when 16#08a5# => read_data_o <= x"3064";
				when 16#08a6# => read_data_o <= x"3064";
				when 16#08a7# => read_data_o <= x"3064";
				when 16#08a8# => read_data_o <= x"3064";
				when 16#08a9# => read_data_o <= x"3064";
				when 16#08aa# => read_data_o <= x"3064";
				when 16#08ab# => read_data_o <= x"3064";
				when 16#08ac# => read_data_o <= x"2000";
				when 16#08ad# => read_data_o <= x"2000";
				when 16#08ae# => read_data_o <= x"2000";
				when 16#08af# => read_data_o <= x"2000";
				when 16#08b0# => read_data_o <= x"2000";
				when 16#08b1# => read_data_o <= x"b196";
				when 16#08b2# => read_data_o <= x"0000";
				when 16#08b3# => read_data_o <= x"0000";
				when 16#08b4# => read_data_o <= x"0000";
				when 16#08b5# => read_data_o <= x"0000";
				when 16#08b6# => read_data_o <= x"0000";
				when 16#08b7# => read_data_o <= x"0000";
				when 16#08b8# => read_data_o <= x"0000";
				when 16#08b9# => read_data_o <= x"0000";
				when 16#08ba# => read_data_o <= x"0000";
				when 16#08bb# => read_data_o <= x"0000";
				when 16#08bc# => read_data_o <= x"0000";
				when 16#08bd# => read_data_o <= x"0000";
				when 16#08be# => read_data_o <= x"0000";
				when 16#08bf# => read_data_o <= x"0000";
				when 16#08c0# => read_data_o <= x"0000";
				when 16#08c1# => read_data_o <= x"0000";
				when 16#08c2# => read_data_o <= x"0000";
				when 16#08c3# => read_data_o <= x"0000";
				when 16#08c4# => read_data_o <= x"0000";
				when 16#08c5# => read_data_o <= x"0000";
				when 16#08c6# => read_data_o <= x"0000";
				when 16#08c7# => read_data_o <= x"0000";
				when 16#08c8# => read_data_o <= x"0000";
				when 16#08c9# => read_data_o <= x"0000";
				when 16#08ca# => read_data_o <= x"0000";
				when 16#08cb# => read_data_o <= x"7064";
				when 16#08cc# => read_data_o <= x"0000";
				when 16#08cd# => read_data_o <= x"0000";
				when 16#08ce# => read_data_o <= x"0000";
				when 16#08cf# => read_data_o <= x"0000";
				when 16#08d0# => read_data_o <= x"0000";
				when 16#08d1# => read_data_o <= x"0000";
				when 16#08d2# => read_data_o <= x"0000";
				when 16#08d3# => read_data_o <= x"0000";
				when 16#08d4# => read_data_o <= x"0000";
				when 16#08d5# => read_data_o <= x"0000";
				when 16#08d6# => read_data_o <= x"0000";
				when 16#08d7# => read_data_o <= x"0000";
				when 16#08d8# => read_data_o <= x"0000";
				when 16#08d9# => read_data_o <= x"0000";
				when 16#08da# => read_data_o <= x"0000";
				when 16#08db# => read_data_o <= x"0000";
				when 16#08dc# => read_data_o <= x"0000";
				when 16#08dd# => read_data_o <= x"0000";
				when 16#08de# => read_data_o <= x"0000";
				when 16#08df# => read_data_o <= x"0000";
				when 16#08e0# => read_data_o <= x"0000";
				when 16#08e1# => read_data_o <= x"0000";
				when 16#08e2# => read_data_o <= x"0000";
				when 16#08e3# => read_data_o <= x"0000";
				when 16#08e4# => read_data_o <= x"0000";
				when 16#08e5# => read_data_o <= x"0000";
				when 16#08e6# => read_data_o <= x"0000";
				when 16#08e7# => read_data_o <= x"0000";
				when 16#08e8# => read_data_o <= x"0000";
				when 16#08e9# => read_data_o <= x"0000";
				when 16#08ea# => read_data_o <= x"0000";
				when 16#08eb# => read_data_o <= x"0000";
				when 16#08ec# => read_data_o <= x"0000";
				when 16#08ed# => read_data_o <= x"0000";
				when 16#08ee# => read_data_o <= x"0000";
				when 16#08ef# => read_data_o <= x"0000";
				when 16#08f0# => read_data_o <= x"0000";
				when 16#08f1# => read_data_o <= x"0000";
				when 16#08f2# => read_data_o <= x"0000";
				when 16#08f3# => read_data_o <= x"0000";
				when 16#08f4# => read_data_o <= x"0000";
				when 16#08f5# => read_data_o <= x"0000";
				when 16#08f6# => read_data_o <= x"0000";
				when 16#08f7# => read_data_o <= x"0000";
				when 16#08f8# => read_data_o <= x"0000";
				when 16#08f9# => read_data_o <= x"0000";
				when 16#08fa# => read_data_o <= x"0000";
				when 16#08fb# => read_data_o <= x"0000";
				when 16#08fc# => read_data_o <= x"0000";
				when 16#08fd# => read_data_o <= x"0000";
				when 16#08fe# => read_data_o <= x"0000";
				when 16#08ff# => read_data_o <= x"0000";
				when 16#0900# => read_data_o <= x"0000";
				when 16#0901# => read_data_o <= x"0000";
				when 16#0902# => read_data_o <= x"0000";
				when 16#0903# => read_data_o <= x"0000";
				when 16#0904# => read_data_o <= x"0000";
				when 16#0905# => read_data_o <= x"0000";
				when 16#0906# => read_data_o <= x"0000";
				when 16#0907# => read_data_o <= x"0000";
				when 16#0908# => read_data_o <= x"0000";
				when 16#0909# => read_data_o <= x"0000";
				when 16#090a# => read_data_o <= x"0000";
				when 16#090b# => read_data_o <= x"0000";
				when 16#090c# => read_data_o <= x"0000";
				when 16#090d# => read_data_o <= x"0000";
				when 16#090e# => read_data_o <= x"0000";
				when 16#090f# => read_data_o <= x"0000";
				when 16#0910# => read_data_o <= x"0000";
				when 16#0911# => read_data_o <= x"0000";
				when 16#0912# => read_data_o <= x"0000";
				when 16#0913# => read_data_o <= x"0000";
				when 16#0914# => read_data_o <= x"0000";
				when 16#0915# => read_data_o <= x"0000";
				when 16#0916# => read_data_o <= x"0000";
				when 16#0917# => read_data_o <= x"0000";
				when 16#0918# => read_data_o <= x"0000";
				when 16#0919# => read_data_o <= x"0000";
				when 16#091a# => read_data_o <= x"0000";
				when 16#091b# => read_data_o <= x"0000";
				when 16#091c# => read_data_o <= x"0000";
				when 16#091d# => read_data_o <= x"0000";
				when 16#091e# => read_data_o <= x"0000";
				when 16#091f# => read_data_o <= x"0000";
				when 16#0920# => read_data_o <= x"0000";
				when 16#0921# => read_data_o <= x"0000";
				when 16#0922# => read_data_o <= x"0000";
				when 16#0923# => read_data_o <= x"0000";
				when 16#0924# => read_data_o <= x"0000";
				when 16#0925# => read_data_o <= x"0000";
				when 16#0926# => read_data_o <= x"0000";
				when 16#0927# => read_data_o <= x"0000";
				when 16#0928# => read_data_o <= x"0000";
				when 16#0929# => read_data_o <= x"0000";
				when 16#092a# => read_data_o <= x"0000";
				when 16#092b# => read_data_o <= x"0000";
				when 16#092c# => read_data_o <= x"0000";
				when 16#092d# => read_data_o <= x"0000";
				when 16#092e# => read_data_o <= x"0000";
				when 16#092f# => read_data_o <= x"0000";
				when 16#0930# => read_data_o <= x"0000";
				when 16#0931# => read_data_o <= x"0000";
				when 16#0932# => read_data_o <= x"0000";
				when 16#0933# => read_data_o <= x"0000";
				when 16#0934# => read_data_o <= x"0000";
				when 16#0935# => read_data_o <= x"0000";
				when 16#0936# => read_data_o <= x"0000";
				when 16#0937# => read_data_o <= x"0000";
				when 16#0938# => read_data_o <= x"0000";
				when 16#0939# => read_data_o <= x"0000";
				when 16#093a# => read_data_o <= x"0000";
				when 16#093b# => read_data_o <= x"0000";
				when 16#093c# => read_data_o <= x"0000";
				when 16#093d# => read_data_o <= x"0000";
				when 16#093e# => read_data_o <= x"0000";
				when 16#093f# => read_data_o <= x"0000";
				when 16#0940# => read_data_o <= x"0000";
				when 16#0941# => read_data_o <= x"0000";
				when 16#0942# => read_data_o <= x"0000";
				when 16#0943# => read_data_o <= x"0000";
				when 16#0944# => read_data_o <= x"0000";
				when 16#0945# => read_data_o <= x"0000";
				when 16#0946# => read_data_o <= x"0000";
				when 16#0947# => read_data_o <= x"0000";
				when 16#0948# => read_data_o <= x"0000";
				when 16#0949# => read_data_o <= x"0000";
				when 16#094a# => read_data_o <= x"0000";
				when 16#094b# => read_data_o <= x"0000";
				when 16#094c# => read_data_o <= x"0000";
				when 16#094d# => read_data_o <= x"0000";
				when 16#094e# => read_data_o <= x"0000";
				when 16#094f# => read_data_o <= x"0000";
				when 16#0950# => read_data_o <= x"0000";
				when 16#0951# => read_data_o <= x"0000";
				when 16#0952# => read_data_o <= x"0000";
				when 16#0953# => read_data_o <= x"0000";
				when 16#0954# => read_data_o <= x"0000";
				when 16#0955# => read_data_o <= x"0000";
				when 16#0956# => read_data_o <= x"0000";
				when 16#0957# => read_data_o <= x"0000";
				when 16#0958# => read_data_o <= x"0000";
				when 16#0959# => read_data_o <= x"0000";
				when 16#095a# => read_data_o <= x"0000";
				when 16#095b# => read_data_o <= x"0000";
				when 16#095c# => read_data_o <= x"0000";
				when 16#095d# => read_data_o <= x"0000";
				when 16#095e# => read_data_o <= x"0000";
				when 16#095f# => read_data_o <= x"0000";
				when 16#0960# => read_data_o <= x"0000";
				when 16#0961# => read_data_o <= x"0000";
				when 16#0962# => read_data_o <= x"0000";
				when 16#0963# => read_data_o <= x"0000";
				when 16#0964# => read_data_o <= x"0000";
				when 16#0965# => read_data_o <= x"0000";
				when 16#0966# => read_data_o <= x"0000";
				when 16#0967# => read_data_o <= x"0000";
				when 16#0968# => read_data_o <= x"0000";
				when 16#0969# => read_data_o <= x"0000";
				when 16#096a# => read_data_o <= x"0000";
				when 16#096b# => read_data_o <= x"0000";
				when 16#096c# => read_data_o <= x"0000";
				when 16#096d# => read_data_o <= x"0000";
				when 16#096e# => read_data_o <= x"0000";
				when 16#096f# => read_data_o <= x"0000";
				when 16#0970# => read_data_o <= x"0000";
				when 16#0971# => read_data_o <= x"0000";
				when 16#0972# => read_data_o <= x"0000";
				when 16#0973# => read_data_o <= x"0000";
				when 16#0974# => read_data_o <= x"0000";
				when 16#0975# => read_data_o <= x"0000";
				when 16#0976# => read_data_o <= x"0000";
				when 16#0977# => read_data_o <= x"0000";
				when 16#0978# => read_data_o <= x"0000";
				when 16#0979# => read_data_o <= x"0000";
				when 16#097a# => read_data_o <= x"0000";
				when 16#097b# => read_data_o <= x"0000";
				when 16#097c# => read_data_o <= x"0000";
				when 16#097d# => read_data_o <= x"0000";
				when 16#097e# => read_data_o <= x"0000";
				when 16#097f# => read_data_o <= x"0000";
				when 16#0980# => read_data_o <= x"0000";
				when 16#0981# => read_data_o <= x"0000";
				when 16#0982# => read_data_o <= x"0000";
				when 16#0983# => read_data_o <= x"0000";
				when 16#0984# => read_data_o <= x"0000";
				when 16#0985# => read_data_o <= x"0000";
				when 16#0986# => read_data_o <= x"0000";
				when 16#0987# => read_data_o <= x"0000";
				when 16#0988# => read_data_o <= x"0000";
				when 16#0989# => read_data_o <= x"0000";
				when 16#098a# => read_data_o <= x"0000";
				when 16#098b# => read_data_o <= x"0000";
				when 16#098c# => read_data_o <= x"0000";
				when 16#098d# => read_data_o <= x"0000";
				when 16#098e# => read_data_o <= x"0000";
				when 16#098f# => read_data_o <= x"0000";
				when 16#0990# => read_data_o <= x"0000";
				when 16#0991# => read_data_o <= x"0000";
				when 16#0992# => read_data_o <= x"0000";
				when 16#0993# => read_data_o <= x"0000";
				when 16#0994# => read_data_o <= x"0000";
				when 16#0995# => read_data_o <= x"0000";
				when 16#0996# => read_data_o <= x"0000";
				when 16#0997# => read_data_o <= x"0000";
				when 16#0998# => read_data_o <= x"0000";
				when 16#0999# => read_data_o <= x"0000";
				when 16#099a# => read_data_o <= x"0000";
				when 16#099b# => read_data_o <= x"0000";
				when 16#099c# => read_data_o <= x"0000";
				when 16#099d# => read_data_o <= x"0000";
				when 16#099e# => read_data_o <= x"0000";
				when 16#099f# => read_data_o <= x"0000";
				when 16#09a0# => read_data_o <= x"0000";
				when 16#09a1# => read_data_o <= x"0000";
				when 16#09a2# => read_data_o <= x"0000";
				when 16#09a3# => read_data_o <= x"0000";
				when 16#09a4# => read_data_o <= x"0000";
				when 16#09a5# => read_data_o <= x"0000";
				when 16#09a6# => read_data_o <= x"0000";
				when 16#09a7# => read_data_o <= x"0000";
				when 16#09a8# => read_data_o <= x"0000";
				when 16#09a9# => read_data_o <= x"0000";
				when 16#09aa# => read_data_o <= x"0000";
				when 16#09ab# => read_data_o <= x"0000";
				when 16#09ac# => read_data_o <= x"0000";
				when 16#09ad# => read_data_o <= x"0000";
				when 16#09ae# => read_data_o <= x"0000";
				when 16#09af# => read_data_o <= x"0000";
				when 16#09b0# => read_data_o <= x"0000";
				when 16#09b1# => read_data_o <= x"0000";
				when 16#09b2# => read_data_o <= x"0000";
				when 16#09b3# => read_data_o <= x"0000";
				when 16#09b4# => read_data_o <= x"0000";
				when 16#09b5# => read_data_o <= x"0000";
				when 16#09b6# => read_data_o <= x"0000";
				when 16#09b7# => read_data_o <= x"0000";
				when 16#09b8# => read_data_o <= x"0000";
				when 16#09b9# => read_data_o <= x"0000";
				when 16#09ba# => read_data_o <= x"0000";
				when 16#09bb# => read_data_o <= x"0000";
				when 16#09bc# => read_data_o <= x"0000";
				when 16#09bd# => read_data_o <= x"0000";
				when 16#09be# => read_data_o <= x"0000";
				when 16#09bf# => read_data_o <= x"0000";
				when 16#09c0# => read_data_o <= x"0000";
				when 16#09c1# => read_data_o <= x"0000";
				when 16#09c2# => read_data_o <= x"0000";
				when 16#09c3# => read_data_o <= x"0000";
				when 16#09c4# => read_data_o <= x"0000";
				when 16#09c5# => read_data_o <= x"0000";
				when 16#09c6# => read_data_o <= x"0000";
				when 16#09c7# => read_data_o <= x"0000";
				when 16#09c8# => read_data_o <= x"0000";
				when 16#09c9# => read_data_o <= x"0000";
				when 16#09ca# => read_data_o <= x"0000";
				when 16#09cb# => read_data_o <= x"0000";
				when 16#09cc# => read_data_o <= x"0000";
				when 16#09cd# => read_data_o <= x"0000";
				when 16#09ce# => read_data_o <= x"0000";
				when 16#09cf# => read_data_o <= x"0000";
				when 16#09d0# => read_data_o <= x"0000";
				when 16#09d1# => read_data_o <= x"0000";
				when 16#09d2# => read_data_o <= x"0000";
				when 16#09d3# => read_data_o <= x"0000";
				when 16#09d4# => read_data_o <= x"0000";
				when 16#09d5# => read_data_o <= x"0000";
				when 16#09d6# => read_data_o <= x"0000";
				when 16#09d7# => read_data_o <= x"0000";
				when 16#09d8# => read_data_o <= x"0000";
				when 16#09d9# => read_data_o <= x"0000";
				when 16#09da# => read_data_o <= x"0000";
				when 16#09db# => read_data_o <= x"0000";
				when 16#09dc# => read_data_o <= x"0000";
				when 16#09dd# => read_data_o <= x"0000";
				when 16#09de# => read_data_o <= x"0000";
				when 16#09df# => read_data_o <= x"0000";
				when 16#09e0# => read_data_o <= x"0000";
				when 16#09e1# => read_data_o <= x"0000";
				when 16#09e2# => read_data_o <= x"0000";
				when 16#09e3# => read_data_o <= x"0000";
				when 16#09e4# => read_data_o <= x"0000";
				when 16#09e5# => read_data_o <= x"0000";
				when 16#09e6# => read_data_o <= x"0000";
				when 16#09e7# => read_data_o <= x"0000";
				when 16#09e8# => read_data_o <= x"0000";
				when 16#09e9# => read_data_o <= x"0000";
				when 16#09ea# => read_data_o <= x"0000";
				when 16#09eb# => read_data_o <= x"0000";
				when 16#09ec# => read_data_o <= x"0000";
				when 16#09ed# => read_data_o <= x"0000";
				when 16#09ee# => read_data_o <= x"0000";
				when 16#09ef# => read_data_o <= x"0000";
				when 16#09f0# => read_data_o <= x"0000";
				when 16#09f1# => read_data_o <= x"0000";
				when 16#09f2# => read_data_o <= x"0000";
				when 16#09f3# => read_data_o <= x"0000";
				when 16#09f4# => read_data_o <= x"0000";
				when 16#09f5# => read_data_o <= x"0000";
				when 16#09f6# => read_data_o <= x"0000";
				when 16#09f7# => read_data_o <= x"0000";
				when 16#09f8# => read_data_o <= x"0000";
				when 16#09f9# => read_data_o <= x"0000";
				when 16#09fa# => read_data_o <= x"0000";
				when 16#09fb# => read_data_o <= x"0000";
				when 16#09fc# => read_data_o <= x"0000";
				when 16#09fd# => read_data_o <= x"0000";
				when 16#09fe# => read_data_o <= x"0000";
				when 16#09ff# => read_data_o <= x"0000";
				when 16#0a00# => read_data_o <= x"0000";
				when 16#0a01# => read_data_o <= x"0000";
				when 16#0a02# => read_data_o <= x"0000";
				when 16#0a03# => read_data_o <= x"0000";
				when 16#0a04# => read_data_o <= x"0000";
				when 16#0a05# => read_data_o <= x"0000";
				when 16#0a06# => read_data_o <= x"0000";
				when 16#0a07# => read_data_o <= x"0000";
				when 16#0a08# => read_data_o <= x"0000";
				when 16#0a09# => read_data_o <= x"0000";
				when 16#0a0a# => read_data_o <= x"0000";
				when 16#0a0b# => read_data_o <= x"0000";
				when 16#0a0c# => read_data_o <= x"0000";
				when 16#0a0d# => read_data_o <= x"0000";
				when 16#0a0e# => read_data_o <= x"0000";
				when 16#0a0f# => read_data_o <= x"0000";
				when 16#0a10# => read_data_o <= x"0000";
				when 16#0a11# => read_data_o <= x"0000";
				when 16#0a12# => read_data_o <= x"0000";
				when 16#0a13# => read_data_o <= x"0000";
				when 16#0a14# => read_data_o <= x"0000";
				when 16#0a15# => read_data_o <= x"0000";
				when 16#0a16# => read_data_o <= x"0000";
				when 16#0a17# => read_data_o <= x"0000";
				when 16#0a18# => read_data_o <= x"0000";
				when 16#0a19# => read_data_o <= x"0000";
				when 16#0a1a# => read_data_o <= x"0000";
				when 16#0a1b# => read_data_o <= x"0000";
				when 16#0a1c# => read_data_o <= x"0000";
				when 16#0a1d# => read_data_o <= x"0000";
				when 16#0a1e# => read_data_o <= x"0000";
				when 16#0a1f# => read_data_o <= x"0000";
				when 16#0a20# => read_data_o <= x"0000";
				when 16#0a21# => read_data_o <= x"0000";
				when 16#0a22# => read_data_o <= x"0000";
				when 16#0a23# => read_data_o <= x"0000";
				when 16#0a24# => read_data_o <= x"0000";
				when 16#0a25# => read_data_o <= x"0000";
				when 16#0a26# => read_data_o <= x"0000";
				when 16#0a27# => read_data_o <= x"0000";
				when 16#0a28# => read_data_o <= x"0000";
				when 16#0a29# => read_data_o <= x"0000";
				when 16#0a2a# => read_data_o <= x"0000";
				when 16#0a2b# => read_data_o <= x"0000";
				when 16#0a2c# => read_data_o <= x"0000";
				when 16#0a2d# => read_data_o <= x"0000";
				when 16#0a2e# => read_data_o <= x"0000";
				when 16#0a2f# => read_data_o <= x"0000";
				when 16#0a30# => read_data_o <= x"0000";
				when 16#0a31# => read_data_o <= x"0000";
				when 16#0a32# => read_data_o <= x"0000";
				when 16#0a33# => read_data_o <= x"0000";
				when 16#0a34# => read_data_o <= x"0000";
				when 16#0a35# => read_data_o <= x"0000";
				when 16#0a36# => read_data_o <= x"0000";
				when 16#0a37# => read_data_o <= x"0000";
				when 16#0a38# => read_data_o <= x"0000";
				when 16#0a39# => read_data_o <= x"0000";
				when 16#0a3a# => read_data_o <= x"0000";
				when 16#0a3b# => read_data_o <= x"0000";
				when 16#0a3c# => read_data_o <= x"0000";
				when 16#0a3d# => read_data_o <= x"0000";
				when 16#0a3e# => read_data_o <= x"0000";
				when 16#0a3f# => read_data_o <= x"0000";
				when 16#0a40# => read_data_o <= x"0000";
				when 16#0a41# => read_data_o <= x"0000";
				when 16#0a42# => read_data_o <= x"0000";
				when 16#0a43# => read_data_o <= x"0000";
				when 16#0a44# => read_data_o <= x"0000";
				when 16#0a45# => read_data_o <= x"0000";
				when 16#0a46# => read_data_o <= x"0000";
				when 16#0a47# => read_data_o <= x"0000";
				when 16#0a48# => read_data_o <= x"0000";
				when 16#0a49# => read_data_o <= x"0000";
				when 16#0a4a# => read_data_o <= x"0000";
				when 16#0a4b# => read_data_o <= x"0000";
				when 16#0a4c# => read_data_o <= x"0000";
				when 16#0a4d# => read_data_o <= x"0000";
				when 16#0a4e# => read_data_o <= x"0000";
				when 16#0a4f# => read_data_o <= x"0000";
				when 16#0a50# => read_data_o <= x"0000";
				when 16#0a51# => read_data_o <= x"0000";
				when 16#0a52# => read_data_o <= x"0000";
				when 16#0a53# => read_data_o <= x"0000";
				when 16#0a54# => read_data_o <= x"0000";
				when 16#0a55# => read_data_o <= x"0000";
				when 16#0a56# => read_data_o <= x"0000";
				when 16#0a57# => read_data_o <= x"0000";
				when 16#0a58# => read_data_o <= x"0000";
				when 16#0a59# => read_data_o <= x"0000";
				when 16#0a5a# => read_data_o <= x"0000";
				when 16#0a5b# => read_data_o <= x"0000";
				when 16#0a5c# => read_data_o <= x"0000";
				when 16#0a5d# => read_data_o <= x"0000";
				when 16#0a5e# => read_data_o <= x"0000";
				when 16#0a5f# => read_data_o <= x"0000";
				when 16#0a60# => read_data_o <= x"0000";
				when 16#0a61# => read_data_o <= x"0000";
				when 16#0a62# => read_data_o <= x"0000";
				when 16#0a63# => read_data_o <= x"0000";
				when 16#0a64# => read_data_o <= x"0000";
				when 16#0a65# => read_data_o <= x"0000";
				when 16#0a66# => read_data_o <= x"0000";
				when 16#0a67# => read_data_o <= x"0000";
				when 16#0a68# => read_data_o <= x"0000";
				when 16#0a69# => read_data_o <= x"0000";
				when 16#0a6a# => read_data_o <= x"0000";
				when 16#0a6b# => read_data_o <= x"0000";
				when 16#0a6c# => read_data_o <= x"0000";
				when 16#0a6d# => read_data_o <= x"0000";
				when 16#0a6e# => read_data_o <= x"0000";
				when 16#0a6f# => read_data_o <= x"0000";
				when 16#0a70# => read_data_o <= x"0000";
				when 16#0a71# => read_data_o <= x"0000";
				when 16#0a72# => read_data_o <= x"0000";
				when 16#0a73# => read_data_o <= x"0000";
				when 16#0a74# => read_data_o <= x"0000";
				when 16#0a75# => read_data_o <= x"0000";
				when 16#0a76# => read_data_o <= x"0000";
				when 16#0a77# => read_data_o <= x"0000";
				when 16#0a78# => read_data_o <= x"0000";
				when 16#0a79# => read_data_o <= x"0000";
				when 16#0a7a# => read_data_o <= x"0000";
				when 16#0a7b# => read_data_o <= x"0000";
				when 16#0a7c# => read_data_o <= x"0000";
				when 16#0a7d# => read_data_o <= x"0000";
				when 16#0a7e# => read_data_o <= x"0000";
				when 16#0a7f# => read_data_o <= x"0000";
				when 16#0a80# => read_data_o <= x"0000";
				when 16#0a81# => read_data_o <= x"0000";
				when 16#0a82# => read_data_o <= x"0000";
				when 16#0a83# => read_data_o <= x"0000";
				when 16#0a84# => read_data_o <= x"0000";
				when 16#0a85# => read_data_o <= x"0000";
				when 16#0a86# => read_data_o <= x"0000";
				when 16#0a87# => read_data_o <= x"0000";
				when 16#0a88# => read_data_o <= x"0000";
				when 16#0a89# => read_data_o <= x"0000";
				when 16#0a8a# => read_data_o <= x"0000";
				when 16#0a8b# => read_data_o <= x"0000";
				when 16#0a8c# => read_data_o <= x"0000";
				when 16#0a8d# => read_data_o <= x"0000";
				when 16#0a8e# => read_data_o <= x"0000";
				when 16#0a8f# => read_data_o <= x"0000";
				when 16#0a90# => read_data_o <= x"0000";
				when 16#0a91# => read_data_o <= x"0000";
				when 16#0a92# => read_data_o <= x"0000";
				when 16#0a93# => read_data_o <= x"0000";
				when 16#0a94# => read_data_o <= x"0000";
				when 16#0a95# => read_data_o <= x"0000";
				when 16#0a96# => read_data_o <= x"0000";
				when 16#0a97# => read_data_o <= x"0000";
				when 16#0a98# => read_data_o <= x"0000";
				when 16#0a99# => read_data_o <= x"0000";
				when 16#0a9a# => read_data_o <= x"0000";
				when 16#0a9b# => read_data_o <= x"0000";
				when 16#0a9c# => read_data_o <= x"0000";
				when 16#0a9d# => read_data_o <= x"0000";
				when 16#0a9e# => read_data_o <= x"0000";
				when 16#0a9f# => read_data_o <= x"0000";
				when 16#0aa0# => read_data_o <= x"0000";
				when 16#0aa1# => read_data_o <= x"0000";
				when 16#0aa2# => read_data_o <= x"0000";
				when 16#0aa3# => read_data_o <= x"0000";
				when 16#0aa4# => read_data_o <= x"0000";
				when 16#0aa5# => read_data_o <= x"0000";
				when 16#0aa6# => read_data_o <= x"0000";
				when 16#0aa7# => read_data_o <= x"0000";
				when 16#0aa8# => read_data_o <= x"0000";
				when 16#0aa9# => read_data_o <= x"0000";
				when 16#0aaa# => read_data_o <= x"0000";
				when 16#0aab# => read_data_o <= x"0000";
				when 16#0aac# => read_data_o <= x"0000";
				when 16#0aad# => read_data_o <= x"0000";
				when 16#0aae# => read_data_o <= x"0000";
				when 16#0aaf# => read_data_o <= x"0000";
				when 16#0ab0# => read_data_o <= x"0000";
				when 16#0ab1# => read_data_o <= x"0000";
				when 16#0ab2# => read_data_o <= x"0000";
				when 16#0ab3# => read_data_o <= x"0000";
				when 16#0ab4# => read_data_o <= x"0000";
				when 16#0ab5# => read_data_o <= x"0000";
				when 16#0ab6# => read_data_o <= x"0000";
				when 16#0ab7# => read_data_o <= x"0000";
				when 16#0ab8# => read_data_o <= x"0000";
				when 16#0ab9# => read_data_o <= x"0000";
				when 16#0aba# => read_data_o <= x"0000";
				when 16#0abb# => read_data_o <= x"0000";
				when 16#0abc# => read_data_o <= x"0000";
				when 16#0abd# => read_data_o <= x"0000";
				when 16#0abe# => read_data_o <= x"0000";
				when 16#0abf# => read_data_o <= x"0000";
				when 16#0ac0# => read_data_o <= x"0000";
				when 16#0ac1# => read_data_o <= x"0000";
				when 16#0ac2# => read_data_o <= x"0000";
				when 16#0ac3# => read_data_o <= x"0000";
				when 16#0ac4# => read_data_o <= x"0000";
				when 16#0ac5# => read_data_o <= x"0000";
				when 16#0ac6# => read_data_o <= x"0000";
				when 16#0ac7# => read_data_o <= x"0000";
				when 16#0ac8# => read_data_o <= x"0000";
				when 16#0ac9# => read_data_o <= x"0000";
				when 16#0aca# => read_data_o <= x"0000";
				when 16#0acb# => read_data_o <= x"0000";
				when 16#0acc# => read_data_o <= x"0000";
				when 16#0acd# => read_data_o <= x"0000";
				when 16#0ace# => read_data_o <= x"0000";
				when 16#0acf# => read_data_o <= x"0000";
				when 16#0ad0# => read_data_o <= x"0000";
				when 16#0ad1# => read_data_o <= x"0000";
				when 16#0ad2# => read_data_o <= x"0000";
				when 16#0ad3# => read_data_o <= x"0000";
				when 16#0ad4# => read_data_o <= x"0000";
				when 16#0ad5# => read_data_o <= x"0000";
				when 16#0ad6# => read_data_o <= x"0000";
				when 16#0ad7# => read_data_o <= x"0000";
				when 16#0ad8# => read_data_o <= x"0000";
				when 16#0ad9# => read_data_o <= x"0000";
				when 16#0ada# => read_data_o <= x"0000";
				when 16#0adb# => read_data_o <= x"0000";
				when 16#0adc# => read_data_o <= x"0000";
				when 16#0add# => read_data_o <= x"0000";
				when 16#0ade# => read_data_o <= x"0000";
				when 16#0adf# => read_data_o <= x"0000";
				when 16#0ae0# => read_data_o <= x"0000";
				when 16#0ae1# => read_data_o <= x"0000";
				when 16#0ae2# => read_data_o <= x"0000";
				when 16#0ae3# => read_data_o <= x"0000";
				when 16#0ae4# => read_data_o <= x"0000";
				when 16#0ae5# => read_data_o <= x"0000";
				when 16#0ae6# => read_data_o <= x"0000";
				when 16#0ae7# => read_data_o <= x"0000";
				when 16#0ae8# => read_data_o <= x"0000";
				when 16#0ae9# => read_data_o <= x"0000";
				when 16#0aea# => read_data_o <= x"0000";
				when 16#0aeb# => read_data_o <= x"0000";
				when 16#0aec# => read_data_o <= x"0000";
				when 16#0aed# => read_data_o <= x"0000";
				when 16#0aee# => read_data_o <= x"0000";
				when 16#0aef# => read_data_o <= x"0000";
				when 16#0af0# => read_data_o <= x"0000";
				when 16#0af1# => read_data_o <= x"0000";
				when 16#0af2# => read_data_o <= x"0000";
				when 16#0af3# => read_data_o <= x"0000";
				when 16#0af4# => read_data_o <= x"0000";
				when 16#0af5# => read_data_o <= x"0000";
				when 16#0af6# => read_data_o <= x"0000";
				when 16#0af7# => read_data_o <= x"0000";
				when 16#0af8# => read_data_o <= x"0000";
				when 16#0af9# => read_data_o <= x"0000";
				when 16#0afa# => read_data_o <= x"0000";
				when 16#0afb# => read_data_o <= x"0000";
				when 16#0afc# => read_data_o <= x"0000";
				when 16#0afd# => read_data_o <= x"0000";
				when 16#0afe# => read_data_o <= x"0000";
				when 16#0aff# => read_data_o <= x"0000";
				when 16#0b00# => read_data_o <= x"0000";
				when 16#0b01# => read_data_o <= x"0000";
				when 16#0b02# => read_data_o <= x"0000";
				when 16#0b03# => read_data_o <= x"0000";
				when 16#0b04# => read_data_o <= x"0000";
				when 16#0b05# => read_data_o <= x"0000";
				when 16#0b06# => read_data_o <= x"0000";
				when 16#0b07# => read_data_o <= x"0000";
				when 16#0b08# => read_data_o <= x"0000";
				when 16#0b09# => read_data_o <= x"0000";
				when 16#0b0a# => read_data_o <= x"0000";
				when 16#0b0b# => read_data_o <= x"0000";
				when 16#0b0c# => read_data_o <= x"0000";
				when 16#0b0d# => read_data_o <= x"0000";
				when 16#0b0e# => read_data_o <= x"0000";
				when 16#0b0f# => read_data_o <= x"0000";
				when 16#0b10# => read_data_o <= x"0000";
				when 16#0b11# => read_data_o <= x"0000";
				when 16#0b12# => read_data_o <= x"0000";
				when 16#0b13# => read_data_o <= x"0000";
				when 16#0b14# => read_data_o <= x"0000";
				when 16#0b15# => read_data_o <= x"0000";
				when 16#0b16# => read_data_o <= x"0000";
				when 16#0b17# => read_data_o <= x"0000";
				when 16#0b18# => read_data_o <= x"0000";
				when 16#0b19# => read_data_o <= x"0000";
				when 16#0b1a# => read_data_o <= x"0000";
				when 16#0b1b# => read_data_o <= x"0000";
				when 16#0b1c# => read_data_o <= x"0000";
				when 16#0b1d# => read_data_o <= x"0000";
				when 16#0b1e# => read_data_o <= x"0000";
				when 16#0b1f# => read_data_o <= x"0000";
				when 16#0b20# => read_data_o <= x"0000";
				when 16#0b21# => read_data_o <= x"0000";
				when 16#0b22# => read_data_o <= x"0000";
				when 16#0b23# => read_data_o <= x"0000";
				when 16#0b24# => read_data_o <= x"0000";
				when 16#0b25# => read_data_o <= x"0000";
				when 16#0b26# => read_data_o <= x"0000";
				when 16#0b27# => read_data_o <= x"0000";
				when 16#0b28# => read_data_o <= x"0000";
				when 16#0b29# => read_data_o <= x"0000";
				when 16#0b2a# => read_data_o <= x"0000";
				when 16#0b2b# => read_data_o <= x"0000";
				when 16#0b2c# => read_data_o <= x"0000";
				when 16#0b2d# => read_data_o <= x"0000";
				when 16#0b2e# => read_data_o <= x"0000";
				when 16#0b2f# => read_data_o <= x"0000";
				when 16#0b30# => read_data_o <= x"0000";
				when 16#0b31# => read_data_o <= x"0000";
				when 16#0b32# => read_data_o <= x"0000";
				when 16#0b33# => read_data_o <= x"0000";
				when 16#0b34# => read_data_o <= x"0000";
				when 16#0b35# => read_data_o <= x"0000";
				when 16#0b36# => read_data_o <= x"0000";
				when 16#0b37# => read_data_o <= x"0000";
				when 16#0b38# => read_data_o <= x"0000";
				when 16#0b39# => read_data_o <= x"0000";
				when 16#0b3a# => read_data_o <= x"0000";
				when 16#0b3b# => read_data_o <= x"0000";
				when 16#0b3c# => read_data_o <= x"0000";
				when 16#0b3d# => read_data_o <= x"0000";
				when 16#0b3e# => read_data_o <= x"0000";
				when 16#0b3f# => read_data_o <= x"0000";
				when 16#0b40# => read_data_o <= x"0000";
				when 16#0b41# => read_data_o <= x"0000";
				when 16#0b42# => read_data_o <= x"0000";
				when 16#0b43# => read_data_o <= x"0000";
				when 16#0b44# => read_data_o <= x"0000";
				when 16#0b45# => read_data_o <= x"0000";
				when 16#0b46# => read_data_o <= x"0000";
				when 16#0b47# => read_data_o <= x"0000";
				when 16#0b48# => read_data_o <= x"0000";
				when 16#0b49# => read_data_o <= x"0000";
				when 16#0b4a# => read_data_o <= x"0000";
				when 16#0b4b# => read_data_o <= x"0000";
				when 16#0b4c# => read_data_o <= x"0000";
				when 16#0b4d# => read_data_o <= x"0000";
				when 16#0b4e# => read_data_o <= x"0000";
				when 16#0b4f# => read_data_o <= x"0000";
				when 16#0b50# => read_data_o <= x"0000";
				when 16#0b51# => read_data_o <= x"0000";
				when 16#0b52# => read_data_o <= x"0000";
				when 16#0b53# => read_data_o <= x"0000";
				when 16#0b54# => read_data_o <= x"0000";
				when 16#0b55# => read_data_o <= x"0000";
				when 16#0b56# => read_data_o <= x"0000";
				when 16#0b57# => read_data_o <= x"0000";
				when 16#0b58# => read_data_o <= x"0000";
				when 16#0b59# => read_data_o <= x"0000";
				when 16#0b5a# => read_data_o <= x"0000";
				when 16#0b5b# => read_data_o <= x"0000";
				when 16#0b5c# => read_data_o <= x"0000";
				when 16#0b5d# => read_data_o <= x"0000";
				when 16#0b5e# => read_data_o <= x"0000";
				when 16#0b5f# => read_data_o <= x"0000";
				when 16#0b60# => read_data_o <= x"0000";
				when 16#0b61# => read_data_o <= x"0000";
				when 16#0b62# => read_data_o <= x"0000";
				when 16#0b63# => read_data_o <= x"0000";
				when 16#0b64# => read_data_o <= x"0000";
				when 16#0b65# => read_data_o <= x"0000";
				when 16#0b66# => read_data_o <= x"0000";
				when 16#0b67# => read_data_o <= x"0000";
				when 16#0b68# => read_data_o <= x"0000";
				when 16#0b69# => read_data_o <= x"0000";
				when 16#0b6a# => read_data_o <= x"0000";
				when 16#0b6b# => read_data_o <= x"0000";
				when 16#0b6c# => read_data_o <= x"0000";
				when 16#0b6d# => read_data_o <= x"0000";
				when 16#0b6e# => read_data_o <= x"0000";
				when 16#0b6f# => read_data_o <= x"0000";
				when 16#0b70# => read_data_o <= x"0000";
				when 16#0b71# => read_data_o <= x"0000";
				when 16#0b72# => read_data_o <= x"0000";
				when 16#0b73# => read_data_o <= x"0000";
				when 16#0b74# => read_data_o <= x"0000";
				when 16#0b75# => read_data_o <= x"0000";
				when 16#0b76# => read_data_o <= x"0000";
				when 16#0b77# => read_data_o <= x"0000";
				when 16#0b78# => read_data_o <= x"0000";
				when 16#0b79# => read_data_o <= x"0000";
				when 16#0b7a# => read_data_o <= x"0000";
				when 16#0b7b# => read_data_o <= x"0000";
				when 16#0b7c# => read_data_o <= x"0000";
				when 16#0b7d# => read_data_o <= x"0000";
				when 16#0b7e# => read_data_o <= x"0000";
				when 16#0b7f# => read_data_o <= x"0000";
				when 16#0b80# => read_data_o <= x"0000";
				when 16#0b81# => read_data_o <= x"0000";
				when 16#0b82# => read_data_o <= x"0000";
				when 16#0b83# => read_data_o <= x"0000";
				when 16#0b84# => read_data_o <= x"0000";
				when 16#0b85# => read_data_o <= x"0000";
				when 16#0b86# => read_data_o <= x"0000";
				when 16#0b87# => read_data_o <= x"0000";
				when 16#0b88# => read_data_o <= x"0000";
				when 16#0b89# => read_data_o <= x"0000";
				when 16#0b8a# => read_data_o <= x"0000";
				when 16#0b8b# => read_data_o <= x"0000";
				when 16#0b8c# => read_data_o <= x"0000";
				when 16#0b8d# => read_data_o <= x"0000";
				when 16#0b8e# => read_data_o <= x"0000";
				when 16#0b8f# => read_data_o <= x"0000";
				when 16#0b90# => read_data_o <= x"0000";
				when 16#0b91# => read_data_o <= x"0000";
				when 16#0b92# => read_data_o <= x"0000";
				when 16#0b93# => read_data_o <= x"0000";
				when 16#0b94# => read_data_o <= x"0000";
				when 16#0b95# => read_data_o <= x"0000";
				when 16#0b96# => read_data_o <= x"0000";
				when 16#0b97# => read_data_o <= x"0000";
				when 16#0b98# => read_data_o <= x"0000";
				when 16#0b99# => read_data_o <= x"0000";
				when 16#0b9a# => read_data_o <= x"0000";
				when 16#0b9b# => read_data_o <= x"0000";
				when 16#0b9c# => read_data_o <= x"0000";
				when 16#0b9d# => read_data_o <= x"0000";
				when 16#0b9e# => read_data_o <= x"0000";
				when 16#0b9f# => read_data_o <= x"0000";
				when 16#0ba0# => read_data_o <= x"0000";
				when 16#0ba1# => read_data_o <= x"0000";
				when 16#0ba2# => read_data_o <= x"0000";
				when 16#0ba3# => read_data_o <= x"0000";
				when 16#0ba4# => read_data_o <= x"0000";
				when 16#0ba5# => read_data_o <= x"0000";
				when 16#0ba6# => read_data_o <= x"0000";
				when 16#0ba7# => read_data_o <= x"0000";
				when 16#0ba8# => read_data_o <= x"0000";
				when 16#0ba9# => read_data_o <= x"0000";
				when 16#0baa# => read_data_o <= x"0000";
				when 16#0bab# => read_data_o <= x"0000";
				when 16#0bac# => read_data_o <= x"0000";
				when 16#0bad# => read_data_o <= x"0000";
				when 16#0bae# => read_data_o <= x"0000";
				when 16#0baf# => read_data_o <= x"0000";
				when 16#0bb0# => read_data_o <= x"0000";
				when 16#0bb1# => read_data_o <= x"0000";
				when 16#0bb2# => read_data_o <= x"0000";
				when 16#0bb3# => read_data_o <= x"0000";
				when 16#0bb4# => read_data_o <= x"0000";
				when 16#0bb5# => read_data_o <= x"0000";
				when 16#0bb6# => read_data_o <= x"0000";
				when 16#0bb7# => read_data_o <= x"0000";
				when 16#0bb8# => read_data_o <= x"0000";
				when 16#0bb9# => read_data_o <= x"0000";
				when 16#0bba# => read_data_o <= x"0000";
				when 16#0bbb# => read_data_o <= x"0000";
				when 16#0bbc# => read_data_o <= x"0000";
				when 16#0bbd# => read_data_o <= x"0000";
				when 16#0bbe# => read_data_o <= x"0000";
				when 16#0bbf# => read_data_o <= x"0000";
				when 16#0bc0# => read_data_o <= x"0000";
				when 16#0bc1# => read_data_o <= x"0000";
				when 16#0bc2# => read_data_o <= x"0000";
				when 16#0bc3# => read_data_o <= x"0000";
				when 16#0bc4# => read_data_o <= x"0000";
				when 16#0bc5# => read_data_o <= x"0000";
				when 16#0bc6# => read_data_o <= x"0000";
				when 16#0bc7# => read_data_o <= x"0000";
				when 16#0bc8# => read_data_o <= x"0000";
				when 16#0bc9# => read_data_o <= x"0000";
				when 16#0bca# => read_data_o <= x"0000";
				when 16#0bcb# => read_data_o <= x"0000";
				when 16#0bcc# => read_data_o <= x"0000";
				when 16#0bcd# => read_data_o <= x"0000";
				when 16#0bce# => read_data_o <= x"0000";
				when 16#0bcf# => read_data_o <= x"0000";
				when 16#0bd0# => read_data_o <= x"0000";
				when 16#0bd1# => read_data_o <= x"0000";
				when 16#0bd2# => read_data_o <= x"0000";
				when 16#0bd3# => read_data_o <= x"0000";
				when 16#0bd4# => read_data_o <= x"0000";
				when 16#0bd5# => read_data_o <= x"0000";
				when 16#0bd6# => read_data_o <= x"0000";
				when 16#0bd7# => read_data_o <= x"0000";
				when 16#0bd8# => read_data_o <= x"0000";
				when 16#0bd9# => read_data_o <= x"0000";
				when 16#0bda# => read_data_o <= x"0000";
				when 16#0bdb# => read_data_o <= x"0000";
				when 16#0bdc# => read_data_o <= x"0000";
				when 16#0bdd# => read_data_o <= x"0000";
				when 16#0bde# => read_data_o <= x"0000";
				when 16#0bdf# => read_data_o <= x"0000";
				when 16#0be0# => read_data_o <= x"0000";
				when 16#0be1# => read_data_o <= x"0000";
				when 16#0be2# => read_data_o <= x"0000";
				when 16#0be3# => read_data_o <= x"0000";
				when 16#0be4# => read_data_o <= x"0000";
				when 16#0be5# => read_data_o <= x"0000";
				when 16#0be6# => read_data_o <= x"0000";
				when 16#0be7# => read_data_o <= x"0000";
				when 16#0be8# => read_data_o <= x"0000";
				when 16#0be9# => read_data_o <= x"0000";
				when 16#0bea# => read_data_o <= x"0000";
				when 16#0beb# => read_data_o <= x"0000";
				when 16#0bec# => read_data_o <= x"0000";
				when 16#0bed# => read_data_o <= x"0000";
				when 16#0bee# => read_data_o <= x"0000";
				when 16#0bef# => read_data_o <= x"0000";
				when 16#0bf0# => read_data_o <= x"0000";
				when 16#0bf1# => read_data_o <= x"0000";
				when 16#0bf2# => read_data_o <= x"0000";
				when 16#0bf3# => read_data_o <= x"0000";
				when 16#0bf4# => read_data_o <= x"0000";
				when 16#0bf5# => read_data_o <= x"0000";
				when 16#0bf6# => read_data_o <= x"0000";
				when 16#0bf7# => read_data_o <= x"0000";
				when 16#0bf8# => read_data_o <= x"0000";
				when 16#0bf9# => read_data_o <= x"0000";
				when 16#0bfa# => read_data_o <= x"0000";
				when 16#0bfb# => read_data_o <= x"0000";
				when 16#0bfc# => read_data_o <= x"0000";
				when 16#0bfd# => read_data_o <= x"0000";
				when 16#0bfe# => read_data_o <= x"0000";
				when 16#0bff# => read_data_o <= x"0000";
				when 16#0c00# => read_data_o <= x"0000";
				when 16#0c01# => read_data_o <= x"0000";
				when 16#0c02# => read_data_o <= x"0000";
				when 16#0c03# => read_data_o <= x"0000";
				when 16#0c04# => read_data_o <= x"0000";
				when 16#0c05# => read_data_o <= x"0000";
				when 16#0c06# => read_data_o <= x"0000";
				when 16#0c07# => read_data_o <= x"0000";
				when 16#0c08# => read_data_o <= x"0000";
				when 16#0c09# => read_data_o <= x"0000";
				when 16#0c0a# => read_data_o <= x"0000";
				when 16#0c0b# => read_data_o <= x"0000";
				when 16#0c0c# => read_data_o <= x"0000";
				when 16#0c0d# => read_data_o <= x"0000";
				when 16#0c0e# => read_data_o <= x"0000";
				when 16#0c0f# => read_data_o <= x"0000";
				when 16#0c10# => read_data_o <= x"0000";
				when 16#0c11# => read_data_o <= x"0000";
				when 16#0c12# => read_data_o <= x"0000";
				when 16#0c13# => read_data_o <= x"0000";
				when 16#0c14# => read_data_o <= x"0000";
				when 16#0c15# => read_data_o <= x"0000";
				when 16#0c16# => read_data_o <= x"0000";
				when 16#0c17# => read_data_o <= x"0000";
				when 16#0c18# => read_data_o <= x"0000";
				when 16#0c19# => read_data_o <= x"0000";
				when 16#0c1a# => read_data_o <= x"0000";
				when 16#0c1b# => read_data_o <= x"0000";
				when 16#0c1c# => read_data_o <= x"0000";
				when 16#0c1d# => read_data_o <= x"0000";
				when 16#0c1e# => read_data_o <= x"0000";
				when 16#0c1f# => read_data_o <= x"0000";
				when 16#0c20# => read_data_o <= x"0000";
				when 16#0c21# => read_data_o <= x"0000";
				when 16#0c22# => read_data_o <= x"0000";
				when 16#0c23# => read_data_o <= x"0000";
				when 16#0c24# => read_data_o <= x"0000";
				when 16#0c25# => read_data_o <= x"0000";
				when 16#0c26# => read_data_o <= x"0000";
				when 16#0c27# => read_data_o <= x"0000";
				when 16#0c28# => read_data_o <= x"0000";
				when 16#0c29# => read_data_o <= x"0000";
				when 16#0c2a# => read_data_o <= x"0000";
				when 16#0c2b# => read_data_o <= x"0000";
				when 16#0c2c# => read_data_o <= x"0000";
				when 16#0c2d# => read_data_o <= x"0000";
				when 16#0c2e# => read_data_o <= x"0000";
				when 16#0c2f# => read_data_o <= x"0000";
				when 16#0c30# => read_data_o <= x"0000";
				when 16#0c31# => read_data_o <= x"0000";
				when 16#0c32# => read_data_o <= x"0000";
				when 16#0c33# => read_data_o <= x"0000";
				when 16#0c34# => read_data_o <= x"0000";
				when 16#0c35# => read_data_o <= x"0000";
				when 16#0c36# => read_data_o <= x"0000";
				when 16#0c37# => read_data_o <= x"0000";
				when 16#0c38# => read_data_o <= x"0000";
				when 16#0c39# => read_data_o <= x"0000";
				when 16#0c3a# => read_data_o <= x"0000";
				when 16#0c3b# => read_data_o <= x"0000";
				when 16#0c3c# => read_data_o <= x"0000";
				when 16#0c3d# => read_data_o <= x"0000";
				when 16#0c3e# => read_data_o <= x"0000";
				when 16#0c3f# => read_data_o <= x"0000";
				when 16#0c40# => read_data_o <= x"0000";
				when 16#0c41# => read_data_o <= x"0000";
				when 16#0c42# => read_data_o <= x"0000";
				when 16#0c43# => read_data_o <= x"0000";
				when 16#0c44# => read_data_o <= x"0000";
				when 16#0c45# => read_data_o <= x"0000";
				when 16#0c46# => read_data_o <= x"0000";
				when 16#0c47# => read_data_o <= x"0000";
				when 16#0c48# => read_data_o <= x"0000";
				when 16#0c49# => read_data_o <= x"0000";
				when 16#0c4a# => read_data_o <= x"0000";
				when 16#0c4b# => read_data_o <= x"0000";
				when 16#0c4c# => read_data_o <= x"0000";
				when 16#0c4d# => read_data_o <= x"0000";
				when 16#0c4e# => read_data_o <= x"0000";
				when 16#0c4f# => read_data_o <= x"0000";
				when 16#0c50# => read_data_o <= x"0000";
				when 16#0c51# => read_data_o <= x"0000";
				when 16#0c52# => read_data_o <= x"0000";
				when 16#0c53# => read_data_o <= x"0000";
				when 16#0c54# => read_data_o <= x"0000";
				when 16#0c55# => read_data_o <= x"0000";
				when 16#0c56# => read_data_o <= x"0000";
				when 16#0c57# => read_data_o <= x"0000";
				when 16#0c58# => read_data_o <= x"0000";
				when 16#0c59# => read_data_o <= x"0000";
				when 16#0c5a# => read_data_o <= x"0000";
				when 16#0c5b# => read_data_o <= x"0000";
				when 16#0c5c# => read_data_o <= x"0000";
				when 16#0c5d# => read_data_o <= x"0000";
				when 16#0c5e# => read_data_o <= x"0000";
				when 16#0c5f# => read_data_o <= x"0000";
				when 16#0c60# => read_data_o <= x"0000";
				when 16#0c61# => read_data_o <= x"0000";
				when 16#0c62# => read_data_o <= x"0000";
				when 16#0c63# => read_data_o <= x"0000";
				when 16#0c64# => read_data_o <= x"0000";
				when 16#0c65# => read_data_o <= x"0000";
				when 16#0c66# => read_data_o <= x"0000";
				when 16#0c67# => read_data_o <= x"0000";
				when 16#0c68# => read_data_o <= x"0000";
				when 16#0c69# => read_data_o <= x"0000";
				when 16#0c6a# => read_data_o <= x"0000";
				when 16#0c6b# => read_data_o <= x"0000";
				when 16#0c6c# => read_data_o <= x"0000";
				when 16#0c6d# => read_data_o <= x"0000";
				when 16#0c6e# => read_data_o <= x"0000";
				when 16#0c6f# => read_data_o <= x"0000";
				when 16#0c70# => read_data_o <= x"0000";
				when 16#0c71# => read_data_o <= x"0000";
				when 16#0c72# => read_data_o <= x"0000";
				when 16#0c73# => read_data_o <= x"0000";
				when 16#0c74# => read_data_o <= x"0000";
				when 16#0c75# => read_data_o <= x"0000";
				when 16#0c76# => read_data_o <= x"0000";
				when 16#0c77# => read_data_o <= x"0000";
				when 16#0c78# => read_data_o <= x"0000";
				when 16#0c79# => read_data_o <= x"0000";
				when 16#0c7a# => read_data_o <= x"0000";
				when 16#0c7b# => read_data_o <= x"0000";
				when 16#0c7c# => read_data_o <= x"0000";
				when 16#0c7d# => read_data_o <= x"0000";
				when 16#0c7e# => read_data_o <= x"0000";
				when 16#0c7f# => read_data_o <= x"0000";
				when 16#0c80# => read_data_o <= x"0000";
				when 16#0c81# => read_data_o <= x"0000";
				when 16#0c82# => read_data_o <= x"0000";
				when 16#0c83# => read_data_o <= x"0000";
				when 16#0c84# => read_data_o <= x"0000";
				when 16#0c85# => read_data_o <= x"0000";
				when 16#0c86# => read_data_o <= x"0000";
				when 16#0c87# => read_data_o <= x"0000";
				when 16#0c88# => read_data_o <= x"0000";
				when 16#0c89# => read_data_o <= x"0000";
				when 16#0c8a# => read_data_o <= x"0000";
				when 16#0c8b# => read_data_o <= x"0000";
				when 16#0c8c# => read_data_o <= x"0000";
				when 16#0c8d# => read_data_o <= x"0000";
				when 16#0c8e# => read_data_o <= x"0000";
				when 16#0c8f# => read_data_o <= x"0000";
				when 16#0c90# => read_data_o <= x"0000";
				when 16#0c91# => read_data_o <= x"0000";
				when 16#0c92# => read_data_o <= x"0000";
				when 16#0c93# => read_data_o <= x"0000";
				when 16#0c94# => read_data_o <= x"0000";
				when 16#0c95# => read_data_o <= x"0000";
				when 16#0c96# => read_data_o <= x"0000";
				when 16#0c97# => read_data_o <= x"0000";
				when 16#0c98# => read_data_o <= x"0000";
				when 16#0c99# => read_data_o <= x"0000";
				when 16#0c9a# => read_data_o <= x"0000";
				when 16#0c9b# => read_data_o <= x"0000";
				when 16#0c9c# => read_data_o <= x"0000";
				when 16#0c9d# => read_data_o <= x"0000";
				when 16#0c9e# => read_data_o <= x"0000";
				when 16#0c9f# => read_data_o <= x"0000";
				when 16#0ca0# => read_data_o <= x"0000";
				when 16#0ca1# => read_data_o <= x"0000";
				when 16#0ca2# => read_data_o <= x"0000";
				when 16#0ca3# => read_data_o <= x"0000";
				when 16#0ca4# => read_data_o <= x"0000";
				when 16#0ca5# => read_data_o <= x"0000";
				when 16#0ca6# => read_data_o <= x"0000";
				when 16#0ca7# => read_data_o <= x"0000";
				when 16#0ca8# => read_data_o <= x"0000";
				when 16#0ca9# => read_data_o <= x"0000";
				when 16#0caa# => read_data_o <= x"0000";
				when 16#0cab# => read_data_o <= x"0000";
				when 16#0cac# => read_data_o <= x"0000";
				when 16#0cad# => read_data_o <= x"0000";
				when 16#0cae# => read_data_o <= x"0000";
				when 16#0caf# => read_data_o <= x"0000";
				when 16#0cb0# => read_data_o <= x"0000";
				when 16#0cb1# => read_data_o <= x"0000";
				when 16#0cb2# => read_data_o <= x"0000";
				when 16#0cb3# => read_data_o <= x"0000";
				when 16#0cb4# => read_data_o <= x"0000";
				when 16#0cb5# => read_data_o <= x"0000";
				when 16#0cb6# => read_data_o <= x"0000";
				when 16#0cb7# => read_data_o <= x"0000";
				when 16#0cb8# => read_data_o <= x"0000";
				when 16#0cb9# => read_data_o <= x"0000";
				when 16#0cba# => read_data_o <= x"0000";
				when 16#0cbb# => read_data_o <= x"0000";
				when 16#0cbc# => read_data_o <= x"0000";
				when 16#0cbd# => read_data_o <= x"0000";
				when 16#0cbe# => read_data_o <= x"0000";
				when 16#0cbf# => read_data_o <= x"0000";
				when 16#0cc0# => read_data_o <= x"0000";
				when 16#0cc1# => read_data_o <= x"0000";
				when 16#0cc2# => read_data_o <= x"0000";
				when 16#0cc3# => read_data_o <= x"0000";
				when 16#0cc4# => read_data_o <= x"0000";
				when 16#0cc5# => read_data_o <= x"0000";
				when 16#0cc6# => read_data_o <= x"0000";
				when 16#0cc7# => read_data_o <= x"0000";
				when 16#0cc8# => read_data_o <= x"0000";
				when 16#0cc9# => read_data_o <= x"0000";
				when 16#0cca# => read_data_o <= x"0000";
				when 16#0ccb# => read_data_o <= x"0000";
				when 16#0ccc# => read_data_o <= x"0000";
				when 16#0ccd# => read_data_o <= x"0000";
				when 16#0cce# => read_data_o <= x"0000";
				when 16#0ccf# => read_data_o <= x"0000";
				when 16#0cd0# => read_data_o <= x"0000";
				when 16#0cd1# => read_data_o <= x"0000";
				when 16#0cd2# => read_data_o <= x"0000";
				when 16#0cd3# => read_data_o <= x"0000";
				when 16#0cd4# => read_data_o <= x"0000";
				when 16#0cd5# => read_data_o <= x"0000";
				when 16#0cd6# => read_data_o <= x"0000";
				when 16#0cd7# => read_data_o <= x"0000";
				when 16#0cd8# => read_data_o <= x"0000";
				when 16#0cd9# => read_data_o <= x"0000";
				when 16#0cda# => read_data_o <= x"0000";
				when 16#0cdb# => read_data_o <= x"0000";
				when 16#0cdc# => read_data_o <= x"0000";
				when 16#0cdd# => read_data_o <= x"0000";
				when 16#0cde# => read_data_o <= x"0000";
				when 16#0cdf# => read_data_o <= x"0000";
				when 16#0ce0# => read_data_o <= x"0000";
				when 16#0ce1# => read_data_o <= x"0000";
				when 16#0ce2# => read_data_o <= x"0000";
				when 16#0ce3# => read_data_o <= x"0000";
				when 16#0ce4# => read_data_o <= x"0000";
				when 16#0ce5# => read_data_o <= x"0000";
				when 16#0ce6# => read_data_o <= x"0000";
				when 16#0ce7# => read_data_o <= x"0000";
				when 16#0ce8# => read_data_o <= x"0000";
				when 16#0ce9# => read_data_o <= x"0000";
				when 16#0cea# => read_data_o <= x"0000";
				when 16#0ceb# => read_data_o <= x"0000";
				when 16#0cec# => read_data_o <= x"0000";
				when 16#0ced# => read_data_o <= x"0000";
				when 16#0cee# => read_data_o <= x"0000";
				when 16#0cef# => read_data_o <= x"0000";
				when 16#0cf0# => read_data_o <= x"0000";
				when 16#0cf1# => read_data_o <= x"0000";
				when 16#0cf2# => read_data_o <= x"0000";
				when 16#0cf3# => read_data_o <= x"0000";
				when 16#0cf4# => read_data_o <= x"0000";
				when 16#0cf5# => read_data_o <= x"0000";
				when 16#0cf6# => read_data_o <= x"0000";
				when 16#0cf7# => read_data_o <= x"0000";
				when 16#0cf8# => read_data_o <= x"0000";
				when 16#0cf9# => read_data_o <= x"0000";
				when 16#0cfa# => read_data_o <= x"0000";
				when 16#0cfb# => read_data_o <= x"0000";
				when 16#0cfc# => read_data_o <= x"0000";
				when 16#0cfd# => read_data_o <= x"0000";
				when 16#0cfe# => read_data_o <= x"0000";
				when 16#0cff# => read_data_o <= x"0000";
				when 16#0d00# => read_data_o <= x"0000";
				when 16#0d01# => read_data_o <= x"0000";
				when 16#0d02# => read_data_o <= x"a000";
				when 16#0d03# => read_data_o <= x"00ec";
				when 16#0d04# => read_data_o <= x"d02b";
				when 16#0d05# => read_data_o <= x"7040";
				when 16#0d06# => read_data_o <= x"00cc";
				when 16#0d07# => read_data_o <= x"d02b";
				when 16#0d08# => read_data_o <= x"7040";
				when 16#0d09# => read_data_o <= x"00ac";
				when 16#0d0a# => read_data_o <= x"d02b";
				when 16#0d0b# => read_data_o <= x"7040";
				when 16#0d0c# => read_data_o <= x"008c";
				when 16#0d0d# => read_data_o <= x"d02b";
				when 16#0d0e# => read_data_o <= x"a4d0";
				when 16#0d0f# => read_data_o <= x"0000";
				when 16#0d10# => read_data_o <= x"0000";
				when 16#0d11# => read_data_o <= x"0000";
				when 16#0d12# => read_data_o <= x"0000";
				when 16#0d13# => read_data_o <= x"0000";
				when 16#0d14# => read_data_o <= x"0000";
				when 16#0d15# => read_data_o <= x"0000";
				when 16#0d16# => read_data_o <= x"0000";
				when 16#0d17# => read_data_o <= x"0000";
				when 16#0d18# => read_data_o <= x"0000";
				when 16#0d19# => read_data_o <= x"0000";
				when 16#0d1a# => read_data_o <= x"0000";
				when 16#0d1b# => read_data_o <= x"0000";
				when 16#0d1c# => read_data_o <= x"0000";
				when 16#0d1d# => read_data_o <= x"0000";
				when 16#0d1e# => read_data_o <= x"0000";
				when 16#0d1f# => read_data_o <= x"0000";
				when 16#0d20# => read_data_o <= x"0000";
				when 16#0d21# => read_data_o <= x"0000";
				when 16#0d22# => read_data_o <= x"0000";
				when 16#0d23# => read_data_o <= x"0000";
				when 16#0d24# => read_data_o <= x"0000";
				when 16#0d25# => read_data_o <= x"0000";
				when 16#0d26# => read_data_o <= x"0000";
				when 16#0d27# => read_data_o <= x"0000";
				when 16#0d28# => read_data_o <= x"0000";
				when 16#0d29# => read_data_o <= x"0000";
				when 16#0d2a# => read_data_o <= x"0000";
				when 16#0d2b# => read_data_o <= x"0000";
				when 16#0d2c# => read_data_o <= x"0000";
				when 16#0d2d# => read_data_o <= x"0000";
				when 16#0d2e# => read_data_o <= x"0000";
				when 16#0d2f# => read_data_o <= x"0000";
				when 16#0d30# => read_data_o <= x"0000";
				when 16#0d31# => read_data_o <= x"0000";
				when 16#0d32# => read_data_o <= x"0000";
				when 16#0d33# => read_data_o <= x"0000";
				when 16#0d34# => read_data_o <= x"0000";
				when 16#0d35# => read_data_o <= x"0000";
				when 16#0d36# => read_data_o <= x"0000";
				when 16#0d37# => read_data_o <= x"0000";
				when 16#0d38# => read_data_o <= x"0000";
				when 16#0d39# => read_data_o <= x"0000";
				when 16#0d3a# => read_data_o <= x"0000";
				when 16#0d3b# => read_data_o <= x"0000";
				when 16#0d3c# => read_data_o <= x"0000";
				when 16#0d3d# => read_data_o <= x"0000";
				when 16#0d3e# => read_data_o <= x"0000";
				when 16#0d3f# => read_data_o <= x"0000";
				when 16#0d40# => read_data_o <= x"0000";
				when 16#0d41# => read_data_o <= x"0000";
				when 16#0d42# => read_data_o <= x"0000";
				when 16#0d43# => read_data_o <= x"0000";
				when 16#0d44# => read_data_o <= x"0000";
				when 16#0d45# => read_data_o <= x"0000";
				when 16#0d46# => read_data_o <= x"0000";
				when 16#0d47# => read_data_o <= x"0000";
				when 16#0d48# => read_data_o <= x"0000";
				when 16#0d49# => read_data_o <= x"0000";
				when 16#0d4a# => read_data_o <= x"0000";
				when 16#0d4b# => read_data_o <= x"0000";
				when 16#0d4c# => read_data_o <= x"0000";
				when 16#0d4d# => read_data_o <= x"0000";
				when 16#0d4e# => read_data_o <= x"0000";
				when 16#0d4f# => read_data_o <= x"0000";
				when 16#0d50# => read_data_o <= x"0000";
				when 16#0d51# => read_data_o <= x"0000";
				when 16#0d52# => read_data_o <= x"0000";
				when 16#0d53# => read_data_o <= x"0000";
				when 16#0d54# => read_data_o <= x"0000";
				when 16#0d55# => read_data_o <= x"0000";
				when 16#0d56# => read_data_o <= x"0000";
				when 16#0d57# => read_data_o <= x"0000";
				when 16#0d58# => read_data_o <= x"0000";
				when 16#0d59# => read_data_o <= x"0000";
				when 16#0d5a# => read_data_o <= x"0000";
				when 16#0d5b# => read_data_o <= x"0000";
				when 16#0d5c# => read_data_o <= x"0000";
				when 16#0d5d# => read_data_o <= x"0000";
				when 16#0d5e# => read_data_o <= x"0000";
				when 16#0d5f# => read_data_o <= x"0000";
				when 16#0d60# => read_data_o <= x"0000";
				when 16#0d61# => read_data_o <= x"0000";
				when 16#0d62# => read_data_o <= x"0000";
				when 16#0d63# => read_data_o <= x"0000";
				when 16#0d64# => read_data_o <= x"0000";
				when 16#0d65# => read_data_o <= x"0000";
				when 16#0d66# => read_data_o <= x"0000";
				when 16#0d67# => read_data_o <= x"0000";
				when 16#0d68# => read_data_o <= x"0000";
				when 16#0d69# => read_data_o <= x"0000";
				when 16#0d6a# => read_data_o <= x"0000";
				when 16#0d6b# => read_data_o <= x"0000";
				when 16#0d6c# => read_data_o <= x"0000";
				when 16#0d6d# => read_data_o <= x"0000";
				when 16#0d6e# => read_data_o <= x"0000";
				when 16#0d6f# => read_data_o <= x"0000";
				when 16#0d70# => read_data_o <= x"0000";
				when 16#0d71# => read_data_o <= x"0000";
				when 16#0d72# => read_data_o <= x"0000";
				when 16#0d73# => read_data_o <= x"0000";
				when 16#0d74# => read_data_o <= x"0000";
				when 16#0d75# => read_data_o <= x"0000";
				when 16#0d76# => read_data_o <= x"0000";
				when 16#0d77# => read_data_o <= x"0000";
				when 16#0d78# => read_data_o <= x"0000";
				when 16#0d79# => read_data_o <= x"0000";
				when 16#0d7a# => read_data_o <= x"0000";
				when 16#0d7b# => read_data_o <= x"0000";
				when 16#0d7c# => read_data_o <= x"0000";
				when 16#0d7d# => read_data_o <= x"0000";
				when 16#0d7e# => read_data_o <= x"0000";
				when 16#0d7f# => read_data_o <= x"0000";
				when 16#0d80# => read_data_o <= x"0000";
				when 16#0d81# => read_data_o <= x"0000";
				when 16#0d82# => read_data_o <= x"0000";
				when 16#0d83# => read_data_o <= x"0000";
				when 16#0d84# => read_data_o <= x"0000";
				when 16#0d85# => read_data_o <= x"0000";
				when 16#0d86# => read_data_o <= x"0000";
				when 16#0d87# => read_data_o <= x"0000";
				when 16#0d88# => read_data_o <= x"0000";
				when 16#0d89# => read_data_o <= x"0000";
				when 16#0d8a# => read_data_o <= x"0000";
				when 16#0d8b# => read_data_o <= x"0000";
				when 16#0d8c# => read_data_o <= x"0000";
				when 16#0d8d# => read_data_o <= x"0000";
				when 16#0d8e# => read_data_o <= x"0000";
				when 16#0d8f# => read_data_o <= x"0000";
				when 16#0d90# => read_data_o <= x"0000";
				when 16#0d91# => read_data_o <= x"0000";
				when 16#0d92# => read_data_o <= x"0000";
				when 16#0d93# => read_data_o <= x"0000";
				when 16#0d94# => read_data_o <= x"0000";
				when 16#0d95# => read_data_o <= x"0000";
				when 16#0d96# => read_data_o <= x"0000";
				when 16#0d97# => read_data_o <= x"0000";
				when 16#0d98# => read_data_o <= x"0000";
				when 16#0d99# => read_data_o <= x"0000";
				when 16#0d9a# => read_data_o <= x"0000";
				when 16#0d9b# => read_data_o <= x"0000";
				when 16#0d9c# => read_data_o <= x"0000";
				when 16#0d9d# => read_data_o <= x"0000";
				when 16#0d9e# => read_data_o <= x"0000";
				when 16#0d9f# => read_data_o <= x"0000";
				when 16#0da0# => read_data_o <= x"0000";
				when 16#0da1# => read_data_o <= x"0000";
				when 16#0da2# => read_data_o <= x"0000";
				when 16#0da3# => read_data_o <= x"0000";
				when 16#0da4# => read_data_o <= x"0000";
				when 16#0da5# => read_data_o <= x"0000";
				when 16#0da6# => read_data_o <= x"0000";
				when 16#0da7# => read_data_o <= x"0000";
				when 16#0da8# => read_data_o <= x"0000";
				when 16#0da9# => read_data_o <= x"0000";
				when 16#0daa# => read_data_o <= x"0000";
				when 16#0dab# => read_data_o <= x"0000";
				when 16#0dac# => read_data_o <= x"0000";
				when 16#0dad# => read_data_o <= x"0000";
				when 16#0dae# => read_data_o <= x"0000";
				when 16#0daf# => read_data_o <= x"0000";
				when 16#0db0# => read_data_o <= x"0000";
				when 16#0db1# => read_data_o <= x"0000";
				when 16#0db2# => read_data_o <= x"0000";
				when 16#0db3# => read_data_o <= x"0000";
				when 16#0db4# => read_data_o <= x"0000";
				when 16#0db5# => read_data_o <= x"0000";
				when 16#0db6# => read_data_o <= x"0000";
				when 16#0db7# => read_data_o <= x"0000";
				when 16#0db8# => read_data_o <= x"0000";
				when 16#0db9# => read_data_o <= x"0000";
				when 16#0dba# => read_data_o <= x"0000";
				when 16#0dbb# => read_data_o <= x"0000";
				when 16#0dbc# => read_data_o <= x"0000";
				when 16#0dbd# => read_data_o <= x"0000";
				when 16#0dbe# => read_data_o <= x"0000";
				when 16#0dbf# => read_data_o <= x"0000";
				when 16#0dc0# => read_data_o <= x"0000";
				when 16#0dc1# => read_data_o <= x"0000";
				when 16#0dc2# => read_data_o <= x"0000";
				when 16#0dc3# => read_data_o <= x"0000";
				when 16#0dc4# => read_data_o <= x"0000";
				when 16#0dc5# => read_data_o <= x"0000";
				when 16#0dc6# => read_data_o <= x"0000";
				when 16#0dc7# => read_data_o <= x"0000";
				when 16#0dc8# => read_data_o <= x"0000";
				when 16#0dc9# => read_data_o <= x"0000";
				when 16#0dca# => read_data_o <= x"0000";
				when 16#0dcb# => read_data_o <= x"0000";
				when 16#0dcc# => read_data_o <= x"0000";
				when 16#0dcd# => read_data_o <= x"0000";
				when 16#0dce# => read_data_o <= x"0000";
				when 16#0dcf# => read_data_o <= x"0000";
				when 16#0dd0# => read_data_o <= x"0000";
				when 16#0dd1# => read_data_o <= x"0000";
				when 16#0dd2# => read_data_o <= x"0000";
				when 16#0dd3# => read_data_o <= x"0000";
				when 16#0dd4# => read_data_o <= x"0000";
				when 16#0dd5# => read_data_o <= x"0000";
				when 16#0dd6# => read_data_o <= x"0000";
				when 16#0dd7# => read_data_o <= x"0000";
				when 16#0dd8# => read_data_o <= x"0000";
				when 16#0dd9# => read_data_o <= x"0000";
				when 16#0dda# => read_data_o <= x"0000";
				when 16#0ddb# => read_data_o <= x"0000";
				when 16#0ddc# => read_data_o <= x"0000";
				when 16#0ddd# => read_data_o <= x"0000";
				when 16#0dde# => read_data_o <= x"0000";
				when 16#0ddf# => read_data_o <= x"0000";
				when 16#0de0# => read_data_o <= x"0000";
				when 16#0de1# => read_data_o <= x"0000";
				when 16#0de2# => read_data_o <= x"0000";
				when 16#0de3# => read_data_o <= x"0000";
				when 16#0de4# => read_data_o <= x"0000";
				when 16#0de5# => read_data_o <= x"0000";
				when 16#0de6# => read_data_o <= x"0000";
				when 16#0de7# => read_data_o <= x"0000";
				when 16#0de8# => read_data_o <= x"0000";
				when 16#0de9# => read_data_o <= x"0000";
				when 16#0dea# => read_data_o <= x"0000";
				when 16#0deb# => read_data_o <= x"0000";
				when 16#0dec# => read_data_o <= x"0000";
				when 16#0ded# => read_data_o <= x"0000";
				when 16#0dee# => read_data_o <= x"0000";
				when 16#0def# => read_data_o <= x"0000";
				when 16#0df0# => read_data_o <= x"0000";
				when 16#0df1# => read_data_o <= x"0000";
				when 16#0df2# => read_data_o <= x"0000";
				when 16#0df3# => read_data_o <= x"0000";
				when 16#0df4# => read_data_o <= x"0000";
				when 16#0df5# => read_data_o <= x"0000";
				when 16#0df6# => read_data_o <= x"0000";
				when 16#0df7# => read_data_o <= x"0000";
				when 16#0df8# => read_data_o <= x"0000";
				when 16#0df9# => read_data_o <= x"0000";
				when 16#0dfa# => read_data_o <= x"0000";
				when 16#0dfb# => read_data_o <= x"0000";
				when 16#0dfc# => read_data_o <= x"0000";
				when 16#0dfd# => read_data_o <= x"0000";
				when 16#0dfe# => read_data_o <= x"0000";
				when 16#0dff# => read_data_o <= x"0000";
				when 16#0e00# => read_data_o <= x"0000";
				when 16#0e01# => read_data_o <= x"0000";
				when 16#0e02# => read_data_o <= x"0000";
				when 16#0e03# => read_data_o <= x"0000";
				when 16#0e04# => read_data_o <= x"0000";
				when 16#0e05# => read_data_o <= x"0000";
				when 16#0e06# => read_data_o <= x"0000";
				when 16#0e07# => read_data_o <= x"0000";
				when 16#0e08# => read_data_o <= x"0000";
				when 16#0e09# => read_data_o <= x"0000";
				when 16#0e0a# => read_data_o <= x"0000";
				when 16#0e0b# => read_data_o <= x"0000";
				when 16#0e0c# => read_data_o <= x"0000";
				when 16#0e0d# => read_data_o <= x"0000";
				when 16#0e0e# => read_data_o <= x"0000";
				when 16#0e0f# => read_data_o <= x"0000";
				when 16#0e10# => read_data_o <= x"0000";
				when 16#0e11# => read_data_o <= x"0000";
				when 16#0e12# => read_data_o <= x"0000";
				when 16#0e13# => read_data_o <= x"0000";
				when 16#0e14# => read_data_o <= x"0000";
				when 16#0e15# => read_data_o <= x"0000";
				when 16#0e16# => read_data_o <= x"0000";
				when 16#0e17# => read_data_o <= x"0000";
				when 16#0e18# => read_data_o <= x"0000";
				when 16#0e19# => read_data_o <= x"0000";
				when 16#0e1a# => read_data_o <= x"0000";
				when 16#0e1b# => read_data_o <= x"0000";
				when 16#0e1c# => read_data_o <= x"0000";
				when 16#0e1d# => read_data_o <= x"0000";
				when 16#0e1e# => read_data_o <= x"0000";
				when 16#0e1f# => read_data_o <= x"0000";
				when 16#0e20# => read_data_o <= x"0000";
				when 16#0e21# => read_data_o <= x"0000";
				when 16#0e22# => read_data_o <= x"0000";
				when 16#0e23# => read_data_o <= x"0000";
				when 16#0e24# => read_data_o <= x"0000";
				when 16#0e25# => read_data_o <= x"0000";
				when 16#0e26# => read_data_o <= x"0000";
				when 16#0e27# => read_data_o <= x"0000";
				when 16#0e28# => read_data_o <= x"0000";
				when 16#0e29# => read_data_o <= x"0000";
				when 16#0e2a# => read_data_o <= x"0000";
				when 16#0e2b# => read_data_o <= x"0000";
				when 16#0e2c# => read_data_o <= x"0000";
				when 16#0e2d# => read_data_o <= x"0000";
				when 16#0e2e# => read_data_o <= x"0000";
				when 16#0e2f# => read_data_o <= x"0000";
				when 16#0e30# => read_data_o <= x"0000";
				when 16#0e31# => read_data_o <= x"0000";
				when 16#0e32# => read_data_o <= x"0000";
				when 16#0e33# => read_data_o <= x"0000";
				when 16#0e34# => read_data_o <= x"0000";
				when 16#0e35# => read_data_o <= x"0000";
				when 16#0e36# => read_data_o <= x"0000";
				when 16#0e37# => read_data_o <= x"0000";
				when 16#0e38# => read_data_o <= x"0000";
				when 16#0e39# => read_data_o <= x"0000";
				when 16#0e3a# => read_data_o <= x"0000";
				when 16#0e3b# => read_data_o <= x"0000";
				when 16#0e3c# => read_data_o <= x"0000";
				when 16#0e3d# => read_data_o <= x"0000";
				when 16#0e3e# => read_data_o <= x"0000";
				when 16#0e3f# => read_data_o <= x"0000";
				when 16#0e40# => read_data_o <= x"0000";
				when 16#0e41# => read_data_o <= x"0000";
				when 16#0e42# => read_data_o <= x"0000";
				when 16#0e43# => read_data_o <= x"0000";
				when 16#0e44# => read_data_o <= x"0000";
				when 16#0e45# => read_data_o <= x"0000";
				when 16#0e46# => read_data_o <= x"0000";
				when 16#0e47# => read_data_o <= x"0000";
				when 16#0e48# => read_data_o <= x"0000";
				when 16#0e49# => read_data_o <= x"0000";
				when 16#0e4a# => read_data_o <= x"0000";
				when 16#0e4b# => read_data_o <= x"0000";
				when 16#0e4c# => read_data_o <= x"0000";
				when 16#0e4d# => read_data_o <= x"0000";
				when 16#0e4e# => read_data_o <= x"0000";
				when 16#0e4f# => read_data_o <= x"0000";
				when 16#0e50# => read_data_o <= x"0000";
				when 16#0e51# => read_data_o <= x"0000";
				when 16#0e52# => read_data_o <= x"0000";
				when 16#0e53# => read_data_o <= x"0000";
				when 16#0e54# => read_data_o <= x"0000";
				when 16#0e55# => read_data_o <= x"0000";
				when 16#0e56# => read_data_o <= x"0000";
				when 16#0e57# => read_data_o <= x"0000";
				when 16#0e58# => read_data_o <= x"0000";
				when 16#0e59# => read_data_o <= x"0000";
				when 16#0e5a# => read_data_o <= x"0000";
				when 16#0e5b# => read_data_o <= x"0000";
				when 16#0e5c# => read_data_o <= x"0000";
				when 16#0e5d# => read_data_o <= x"0000";
				when 16#0e5e# => read_data_o <= x"0000";
				when 16#0e5f# => read_data_o <= x"0000";
				when 16#0e60# => read_data_o <= x"0000";
				when 16#0e61# => read_data_o <= x"0000";
				when 16#0e62# => read_data_o <= x"0000";
				when 16#0e63# => read_data_o <= x"0000";
				when 16#0e64# => read_data_o <= x"0000";
				when 16#0e65# => read_data_o <= x"0000";
				when 16#0e66# => read_data_o <= x"0000";
				when 16#0e67# => read_data_o <= x"0000";
				when 16#0e68# => read_data_o <= x"0000";
				when 16#0e69# => read_data_o <= x"0000";
				when 16#0e6a# => read_data_o <= x"0000";
				when 16#0e6b# => read_data_o <= x"0000";
				when 16#0e6c# => read_data_o <= x"0000";
				when 16#0e6d# => read_data_o <= x"0000";
				when 16#0e6e# => read_data_o <= x"0000";
				when 16#0e6f# => read_data_o <= x"0000";
				when 16#0e70# => read_data_o <= x"0000";
				when 16#0e71# => read_data_o <= x"0000";
				when 16#0e72# => read_data_o <= x"0000";
				when 16#0e73# => read_data_o <= x"0000";
				when 16#0e74# => read_data_o <= x"0000";
				when 16#0e75# => read_data_o <= x"0000";
				when 16#0e76# => read_data_o <= x"0000";
				when 16#0e77# => read_data_o <= x"0000";
				when 16#0e78# => read_data_o <= x"0000";
				when 16#0e79# => read_data_o <= x"0000";
				when 16#0e7a# => read_data_o <= x"0000";
				when 16#0e7b# => read_data_o <= x"0000";
				when 16#0e7c# => read_data_o <= x"0000";
				when 16#0e7d# => read_data_o <= x"0000";
				when 16#0e7e# => read_data_o <= x"0000";
				when 16#0e7f# => read_data_o <= x"0000";
				when 16#0e80# => read_data_o <= x"0000";
				when 16#0e81# => read_data_o <= x"0000";
				when 16#0e82# => read_data_o <= x"0000";
				when 16#0e83# => read_data_o <= x"0000";
				when 16#0e84# => read_data_o <= x"0000";
				when 16#0e85# => read_data_o <= x"0000";
				when 16#0e86# => read_data_o <= x"0000";
				when 16#0e87# => read_data_o <= x"0000";
				when 16#0e88# => read_data_o <= x"0000";
				when 16#0e89# => read_data_o <= x"0000";
				when 16#0e8a# => read_data_o <= x"0000";
				when 16#0e8b# => read_data_o <= x"0000";
				when 16#0e8c# => read_data_o <= x"0000";
				when 16#0e8d# => read_data_o <= x"0000";
				when 16#0e8e# => read_data_o <= x"0000";
				when 16#0e8f# => read_data_o <= x"0000";
				when 16#0e90# => read_data_o <= x"0000";
				when 16#0e91# => read_data_o <= x"0000";
				when 16#0e92# => read_data_o <= x"0000";
				when 16#0e93# => read_data_o <= x"0000";
				when 16#0e94# => read_data_o <= x"0000";
				when 16#0e95# => read_data_o <= x"0000";
				when 16#0e96# => read_data_o <= x"0000";
				when 16#0e97# => read_data_o <= x"0000";
				when 16#0e98# => read_data_o <= x"0000";
				when 16#0e99# => read_data_o <= x"0000";
				when 16#0e9a# => read_data_o <= x"0000";
				when 16#0e9b# => read_data_o <= x"0000";
				when 16#0e9c# => read_data_o <= x"0000";
				when 16#0e9d# => read_data_o <= x"0000";
				when 16#0e9e# => read_data_o <= x"0000";
				when 16#0e9f# => read_data_o <= x"0000";
				when 16#0ea0# => read_data_o <= x"0000";
				when 16#0ea1# => read_data_o <= x"0000";
				when 16#0ea2# => read_data_o <= x"0000";
				when 16#0ea3# => read_data_o <= x"0000";
				when 16#0ea4# => read_data_o <= x"0000";
				when 16#0ea5# => read_data_o <= x"0000";
				when 16#0ea6# => read_data_o <= x"0000";
				when 16#0ea7# => read_data_o <= x"0000";
				when 16#0ea8# => read_data_o <= x"0000";
				when 16#0ea9# => read_data_o <= x"0000";
				when 16#0eaa# => read_data_o <= x"0000";
				when 16#0eab# => read_data_o <= x"0000";
				when 16#0eac# => read_data_o <= x"0000";
				when 16#0ead# => read_data_o <= x"0000";
				when 16#0eae# => read_data_o <= x"0000";
				when 16#0eaf# => read_data_o <= x"0000";
				when 16#0eb0# => read_data_o <= x"0000";
				when 16#0eb1# => read_data_o <= x"0000";
				when 16#0eb2# => read_data_o <= x"0000";
				when 16#0eb3# => read_data_o <= x"0000";
				when 16#0eb4# => read_data_o <= x"0000";
				when 16#0eb5# => read_data_o <= x"0000";
				when 16#0eb6# => read_data_o <= x"0000";
				when 16#0eb7# => read_data_o <= x"0000";
				when 16#0eb8# => read_data_o <= x"0000";
				when 16#0eb9# => read_data_o <= x"0000";
				when 16#0eba# => read_data_o <= x"0000";
				when 16#0ebb# => read_data_o <= x"0000";
				when 16#0ebc# => read_data_o <= x"0000";
				when 16#0ebd# => read_data_o <= x"0000";
				when 16#0ebe# => read_data_o <= x"0000";
				when 16#0ebf# => read_data_o <= x"0000";
				when 16#0ec0# => read_data_o <= x"0000";
				when 16#0ec1# => read_data_o <= x"0000";
				when 16#0ec2# => read_data_o <= x"0000";
				when 16#0ec3# => read_data_o <= x"0000";
				when 16#0ec4# => read_data_o <= x"0000";
				when 16#0ec5# => read_data_o <= x"0000";
				when 16#0ec6# => read_data_o <= x"0000";
				when 16#0ec7# => read_data_o <= x"0000";
				when 16#0ec8# => read_data_o <= x"0000";
				when 16#0ec9# => read_data_o <= x"0000";
				when 16#0eca# => read_data_o <= x"0000";
				when 16#0ecb# => read_data_o <= x"0000";
				when 16#0ecc# => read_data_o <= x"0000";
				when 16#0ecd# => read_data_o <= x"0000";
				when 16#0ece# => read_data_o <= x"0000";
				when 16#0ecf# => read_data_o <= x"0000";
				when 16#0ed0# => read_data_o <= x"0000";
				when 16#0ed1# => read_data_o <= x"0000";
				when 16#0ed2# => read_data_o <= x"0000";
				when 16#0ed3# => read_data_o <= x"0000";
				when 16#0ed4# => read_data_o <= x"0000";
				when 16#0ed5# => read_data_o <= x"0000";
				when 16#0ed6# => read_data_o <= x"0000";
				when 16#0ed7# => read_data_o <= x"0000";
				when 16#0ed8# => read_data_o <= x"0000";
				when 16#0ed9# => read_data_o <= x"0000";
				when 16#0eda# => read_data_o <= x"0000";
				when 16#0edb# => read_data_o <= x"0000";
				when 16#0edc# => read_data_o <= x"0000";
				when 16#0edd# => read_data_o <= x"0000";
				when 16#0ede# => read_data_o <= x"0000";
				when 16#0edf# => read_data_o <= x"0000";
				when 16#0ee0# => read_data_o <= x"0000";
				when 16#0ee1# => read_data_o <= x"0000";
				when 16#0ee2# => read_data_o <= x"0000";
				when 16#0ee3# => read_data_o <= x"0000";
				when 16#0ee4# => read_data_o <= x"0000";
				when 16#0ee5# => read_data_o <= x"0000";
				when 16#0ee6# => read_data_o <= x"0000";
				when 16#0ee7# => read_data_o <= x"0000";
				when 16#0ee8# => read_data_o <= x"0000";
				when 16#0ee9# => read_data_o <= x"0000";
				when 16#0eea# => read_data_o <= x"0000";
				when 16#0eeb# => read_data_o <= x"0000";
				when 16#0eec# => read_data_o <= x"0000";
				when 16#0eed# => read_data_o <= x"0000";
				when 16#0eee# => read_data_o <= x"0000";
				when 16#0eef# => read_data_o <= x"0000";
				when 16#0ef0# => read_data_o <= x"0000";
				when 16#0ef1# => read_data_o <= x"0000";
				when 16#0ef2# => read_data_o <= x"0000";
				when 16#0ef3# => read_data_o <= x"0000";
				when 16#0ef4# => read_data_o <= x"0000";
				when 16#0ef5# => read_data_o <= x"0000";
				when 16#0ef6# => read_data_o <= x"0000";
				when 16#0ef7# => read_data_o <= x"0000";
				when 16#0ef8# => read_data_o <= x"0000";
				when 16#0ef9# => read_data_o <= x"0000";
				when 16#0efa# => read_data_o <= x"0000";
				when 16#0efb# => read_data_o <= x"0000";
				when 16#0efc# => read_data_o <= x"0000";
				when 16#0efd# => read_data_o <= x"0000";
				when 16#0efe# => read_data_o <= x"0000";
				when 16#0eff# => read_data_o <= x"0000";
				when 16#0f00# => read_data_o <= x"0000";
				when 16#0f01# => read_data_o <= x"0000";
				when 16#0f02# => read_data_o <= x"0000";
				when 16#0f03# => read_data_o <= x"0000";
				when 16#0f04# => read_data_o <= x"0000";
				when 16#0f05# => read_data_o <= x"0000";
				when 16#0f06# => read_data_o <= x"0000";
				when 16#0f07# => read_data_o <= x"0000";
				when 16#0f08# => read_data_o <= x"0000";
				when 16#0f09# => read_data_o <= x"0000";
				when 16#0f0a# => read_data_o <= x"0000";
				when 16#0f0b# => read_data_o <= x"0000";
				when 16#0f0c# => read_data_o <= x"0000";
				when 16#0f0d# => read_data_o <= x"0000";
				when 16#0f0e# => read_data_o <= x"0000";
				when 16#0f0f# => read_data_o <= x"0000";
				when 16#0f10# => read_data_o <= x"0000";
				when 16#0f11# => read_data_o <= x"0000";
				when 16#0f12# => read_data_o <= x"0000";
				when 16#0f13# => read_data_o <= x"0000";
				when 16#0f14# => read_data_o <= x"0000";
				when 16#0f15# => read_data_o <= x"0000";
				when 16#0f16# => read_data_o <= x"0000";
				when 16#0f17# => read_data_o <= x"0000";
				when 16#0f18# => read_data_o <= x"0000";
				when 16#0f19# => read_data_o <= x"0000";
				when 16#0f1a# => read_data_o <= x"0000";
				when 16#0f1b# => read_data_o <= x"0000";
				when 16#0f1c# => read_data_o <= x"0000";
				when 16#0f1d# => read_data_o <= x"0000";
				when 16#0f1e# => read_data_o <= x"0000";
				when 16#0f1f# => read_data_o <= x"0000";
				when 16#0f20# => read_data_o <= x"0000";
				when 16#0f21# => read_data_o <= x"0000";
				when 16#0f22# => read_data_o <= x"0000";
				when 16#0f23# => read_data_o <= x"0000";
				when 16#0f24# => read_data_o <= x"0000";
				when 16#0f25# => read_data_o <= x"0000";
				when 16#0f26# => read_data_o <= x"0000";
				when 16#0f27# => read_data_o <= x"0000";
				when 16#0f28# => read_data_o <= x"0000";
				when 16#0f29# => read_data_o <= x"0000";
				when 16#0f2a# => read_data_o <= x"0000";
				when 16#0f2b# => read_data_o <= x"0000";
				when 16#0f2c# => read_data_o <= x"0000";
				when 16#0f2d# => read_data_o <= x"0000";
				when 16#0f2e# => read_data_o <= x"0000";
				when 16#0f2f# => read_data_o <= x"0000";
				when 16#0f30# => read_data_o <= x"0000";
				when 16#0f31# => read_data_o <= x"0000";
				when 16#0f32# => read_data_o <= x"0000";
				when 16#0f33# => read_data_o <= x"0000";
				when 16#0f34# => read_data_o <= x"0000";
				when 16#0f35# => read_data_o <= x"0000";
				when 16#0f36# => read_data_o <= x"0000";
				when 16#0f37# => read_data_o <= x"0000";
				when 16#0f38# => read_data_o <= x"0000";
				when 16#0f39# => read_data_o <= x"0000";
				when 16#0f3a# => read_data_o <= x"0000";
				when 16#0f3b# => read_data_o <= x"0000";
				when 16#0f3c# => read_data_o <= x"0000";
				when 16#0f3d# => read_data_o <= x"0000";
				when 16#0f3e# => read_data_o <= x"0000";
				when 16#0f3f# => read_data_o <= x"0000";
				when 16#0f40# => read_data_o <= x"0000";
				when 16#0f41# => read_data_o <= x"0000";
				when 16#0f42# => read_data_o <= x"0000";
				when 16#0f43# => read_data_o <= x"0000";
				when 16#0f44# => read_data_o <= x"0000";
				when 16#0f45# => read_data_o <= x"0000";
				when 16#0f46# => read_data_o <= x"0000";
				when 16#0f47# => read_data_o <= x"0000";
				when 16#0f48# => read_data_o <= x"0000";
				when 16#0f49# => read_data_o <= x"0000";
				when 16#0f4a# => read_data_o <= x"0000";
				when 16#0f4b# => read_data_o <= x"0000";
				when 16#0f4c# => read_data_o <= x"0000";
				when 16#0f4d# => read_data_o <= x"0000";
				when 16#0f4e# => read_data_o <= x"0000";
				when 16#0f4f# => read_data_o <= x"0000";
				when 16#0f50# => read_data_o <= x"0000";
				when 16#0f51# => read_data_o <= x"0000";
				when 16#0f52# => read_data_o <= x"0000";
				when 16#0f53# => read_data_o <= x"0000";
				when 16#0f54# => read_data_o <= x"0000";
				when 16#0f55# => read_data_o <= x"0000";
				when 16#0f56# => read_data_o <= x"0000";
				when 16#0f57# => read_data_o <= x"0000";
				when 16#0f58# => read_data_o <= x"0000";
				when 16#0f59# => read_data_o <= x"0000";
				when 16#0f5a# => read_data_o <= x"0000";
				when 16#0f5b# => read_data_o <= x"0000";
				when 16#0f5c# => read_data_o <= x"0000";
				when 16#0f5d# => read_data_o <= x"0000";
				when 16#0f5e# => read_data_o <= x"0000";
				when 16#0f5f# => read_data_o <= x"0000";
				when 16#0f60# => read_data_o <= x"0000";
				when 16#0f61# => read_data_o <= x"0000";
				when 16#0f62# => read_data_o <= x"0000";
				when 16#0f63# => read_data_o <= x"0000";
				when 16#0f64# => read_data_o <= x"0000";
				when 16#0f65# => read_data_o <= x"0000";
				when 16#0f66# => read_data_o <= x"0000";
				when 16#0f67# => read_data_o <= x"0000";
				when 16#0f68# => read_data_o <= x"0000";
				when 16#0f69# => read_data_o <= x"0000";
				when 16#0f6a# => read_data_o <= x"0000";
				when 16#0f6b# => read_data_o <= x"0000";
				when 16#0f6c# => read_data_o <= x"0000";
				when 16#0f6d# => read_data_o <= x"0000";
				when 16#0f6e# => read_data_o <= x"0000";
				when 16#0f6f# => read_data_o <= x"0000";
				when 16#0f70# => read_data_o <= x"0000";
				when 16#0f71# => read_data_o <= x"0000";
				when 16#0f72# => read_data_o <= x"0000";
				when 16#0f73# => read_data_o <= x"0000";
				when 16#0f74# => read_data_o <= x"0000";
				when 16#0f75# => read_data_o <= x"0000";
				when 16#0f76# => read_data_o <= x"0000";
				when 16#0f77# => read_data_o <= x"0000";
				when 16#0f78# => read_data_o <= x"0000";
				when 16#0f79# => read_data_o <= x"0000";
				when 16#0f7a# => read_data_o <= x"0000";
				when 16#0f7b# => read_data_o <= x"0000";
				when 16#0f7c# => read_data_o <= x"0000";
				when 16#0f7d# => read_data_o <= x"0000";
				when 16#0f7e# => read_data_o <= x"0000";
				when 16#0f7f# => read_data_o <= x"0000";
				when 16#0f80# => read_data_o <= x"0000";
				when 16#0f81# => read_data_o <= x"0000";
				when 16#0f82# => read_data_o <= x"0000";
				when 16#0f83# => read_data_o <= x"0000";
				when 16#0f84# => read_data_o <= x"0000";
				when 16#0f85# => read_data_o <= x"0000";
				when 16#0f86# => read_data_o <= x"0000";
				when 16#0f87# => read_data_o <= x"0000";
				when 16#0f88# => read_data_o <= x"0000";
				when 16#0f89# => read_data_o <= x"0000";
				when 16#0f8a# => read_data_o <= x"0000";
				when 16#0f8b# => read_data_o <= x"0000";
				when 16#0f8c# => read_data_o <= x"0000";
				when 16#0f8d# => read_data_o <= x"0000";
				when 16#0f8e# => read_data_o <= x"0000";
				when 16#0f8f# => read_data_o <= x"0000";
				when 16#0f90# => read_data_o <= x"0000";
				when 16#0f91# => read_data_o <= x"0000";
				when 16#0f92# => read_data_o <= x"0000";
				when 16#0f93# => read_data_o <= x"0000";
				when 16#0f94# => read_data_o <= x"0000";
				when 16#0f95# => read_data_o <= x"0000";
				when 16#0f96# => read_data_o <= x"0000";
				when 16#0f97# => read_data_o <= x"0000";
				when 16#0f98# => read_data_o <= x"0000";
				when 16#0f99# => read_data_o <= x"0000";
				when 16#0f9a# => read_data_o <= x"0000";
				when 16#0f9b# => read_data_o <= x"0000";
				when 16#0f9c# => read_data_o <= x"0000";
				when 16#0f9d# => read_data_o <= x"0000";
				when 16#0f9e# => read_data_o <= x"0000";
				when 16#0f9f# => read_data_o <= x"0000";
				when 16#0fa0# => read_data_o <= x"0000";
				when 16#0fa1# => read_data_o <= x"0000";
				when 16#0fa2# => read_data_o <= x"0000";
				when 16#0fa3# => read_data_o <= x"0000";
				when 16#0fa4# => read_data_o <= x"0000";
				when 16#0fa5# => read_data_o <= x"0000";
				when 16#0fa6# => read_data_o <= x"0000";
				when 16#0fa7# => read_data_o <= x"0000";
				when 16#0fa8# => read_data_o <= x"0000";
				when 16#0fa9# => read_data_o <= x"0000";
				when 16#0faa# => read_data_o <= x"0000";
				when 16#0fab# => read_data_o <= x"0000";
				when 16#0fac# => read_data_o <= x"0000";
				when 16#0fad# => read_data_o <= x"0000";
				when 16#0fae# => read_data_o <= x"0000";
				when 16#0faf# => read_data_o <= x"0000";
				when 16#0fb0# => read_data_o <= x"0000";
				when 16#0fb1# => read_data_o <= x"0000";
				when 16#0fb2# => read_data_o <= x"0000";
				when 16#0fb3# => read_data_o <= x"0000";
				when 16#0fb4# => read_data_o <= x"0000";
				when 16#0fb5# => read_data_o <= x"0000";
				when 16#0fb6# => read_data_o <= x"0000";
				when 16#0fb7# => read_data_o <= x"0000";
				when 16#0fb8# => read_data_o <= x"0000";
				when 16#0fb9# => read_data_o <= x"0000";
				when 16#0fba# => read_data_o <= x"0000";
				when 16#0fbb# => read_data_o <= x"0000";
				when 16#0fbc# => read_data_o <= x"0000";
				when 16#0fbd# => read_data_o <= x"0000";
				when 16#0fbe# => read_data_o <= x"0000";
				when 16#0fbf# => read_data_o <= x"0000";
				when 16#0fc0# => read_data_o <= x"0000";
				when 16#0fc1# => read_data_o <= x"0000";
				when 16#0fc2# => read_data_o <= x"0000";
				when 16#0fc3# => read_data_o <= x"0000";
				when 16#0fc4# => read_data_o <= x"0000";
				when 16#0fc5# => read_data_o <= x"0000";
				when 16#0fc6# => read_data_o <= x"0000";
				when 16#0fc7# => read_data_o <= x"0000";
				when 16#0fc8# => read_data_o <= x"0000";
				when 16#0fc9# => read_data_o <= x"0000";
				when 16#0fca# => read_data_o <= x"0000";
				when 16#0fcb# => read_data_o <= x"0000";
				when 16#0fcc# => read_data_o <= x"0000";
				when 16#0fcd# => read_data_o <= x"0000";
				when 16#0fce# => read_data_o <= x"0000";
				when 16#0fcf# => read_data_o <= x"0000";
				when 16#0fd0# => read_data_o <= x"0000";
				when 16#0fd1# => read_data_o <= x"0000";
				when 16#0fd2# => read_data_o <= x"0000";
				when 16#0fd3# => read_data_o <= x"0000";
				when 16#0fd4# => read_data_o <= x"0000";
				when 16#0fd5# => read_data_o <= x"0000";
				when 16#0fd6# => read_data_o <= x"0000";
				when 16#0fd7# => read_data_o <= x"0000";
				when 16#0fd8# => read_data_o <= x"0000";
				when 16#0fd9# => read_data_o <= x"0000";
				when 16#0fda# => read_data_o <= x"0000";
				when 16#0fdb# => read_data_o <= x"0000";
				when 16#0fdc# => read_data_o <= x"0000";
				when 16#0fdd# => read_data_o <= x"0000";
				when 16#0fde# => read_data_o <= x"0000";
				when 16#0fdf# => read_data_o <= x"0000";
				when 16#0fe0# => read_data_o <= x"0000";
				when 16#0fe1# => read_data_o <= x"0000";
				when 16#0fe2# => read_data_o <= x"0000";
				when 16#0fe3# => read_data_o <= x"0000";
				when 16#0fe4# => read_data_o <= x"0000";
				when 16#0fe5# => read_data_o <= x"0000";
				when 16#0fe6# => read_data_o <= x"0000";
				when 16#0fe7# => read_data_o <= x"0000";
				when 16#0fe8# => read_data_o <= x"0000";
				when 16#0fe9# => read_data_o <= x"0000";
				when 16#0fea# => read_data_o <= x"0000";
				when 16#0feb# => read_data_o <= x"0000";
				when 16#0fec# => read_data_o <= x"0000";
				when 16#0fed# => read_data_o <= x"0000";
				when 16#0fee# => read_data_o <= x"0000";
				when 16#0fef# => read_data_o <= x"0000";
				when 16#0ff0# => read_data_o <= x"0000";
				when 16#0ff1# => read_data_o <= x"0000";
				when 16#0ff2# => read_data_o <= x"0000";
				when 16#0ff3# => read_data_o <= x"0000";
				when 16#0ff4# => read_data_o <= x"0000";
				when 16#0ff5# => read_data_o <= x"0000";
				when 16#0ff6# => read_data_o <= x"0000";
				when 16#0ff7# => read_data_o <= x"0000";
				when 16#0ff8# => read_data_o <= x"0000";
				when 16#0ff9# => read_data_o <= x"0000";
				when 16#0ffa# => read_data_o <= x"0000";
				when 16#0ffb# => read_data_o <= x"0000";
				when 16#0ffc# => read_data_o <= x"0000";
				when 16#0ffd# => read_data_o <= x"0000";
				when 16#0ffe# => read_data_o <= x"0000";
				when 16#0fff# => read_data_o <= x"0000";
				when 16#1000# => read_data_o <= x"0000";
				when 16#1001# => read_data_o <= x"0000";
				when 16#1002# => read_data_o <= x"0000";
				when 16#1003# => read_data_o <= x"0000";
				when 16#1004# => read_data_o <= x"0000";
				when 16#1005# => read_data_o <= x"0000";
				when 16#1006# => read_data_o <= x"0000";
				when 16#1007# => read_data_o <= x"0000";
				when 16#1008# => read_data_o <= x"0000";
				when 16#1009# => read_data_o <= x"0000";
				when 16#100a# => read_data_o <= x"0000";
				when 16#100b# => read_data_o <= x"0000";
				when 16#100c# => read_data_o <= x"0000";
				when 16#100d# => read_data_o <= x"0000";
				when 16#100e# => read_data_o <= x"0000";
				when 16#100f# => read_data_o <= x"0000";
				when 16#1010# => read_data_o <= x"0000";
				when 16#1011# => read_data_o <= x"0000";
				when 16#1012# => read_data_o <= x"0000";
				when 16#1013# => read_data_o <= x"0000";
				when 16#1014# => read_data_o <= x"0000";
				when 16#1015# => read_data_o <= x"0000";
				when 16#1016# => read_data_o <= x"0000";
				when 16#1017# => read_data_o <= x"0000";
				when 16#1018# => read_data_o <= x"0000";
				when 16#1019# => read_data_o <= x"0000";
				when 16#101a# => read_data_o <= x"0000";
				when 16#101b# => read_data_o <= x"0000";
				when 16#101c# => read_data_o <= x"0000";
				when 16#101d# => read_data_o <= x"0000";
				when 16#101e# => read_data_o <= x"0000";
				when 16#101f# => read_data_o <= x"0000";
				when 16#1020# => read_data_o <= x"0000";
				when 16#1021# => read_data_o <= x"0000";
				when 16#1022# => read_data_o <= x"0000";
				when 16#1023# => read_data_o <= x"0000";
				when 16#1024# => read_data_o <= x"0000";
				when 16#1025# => read_data_o <= x"0000";
				when 16#1026# => read_data_o <= x"0000";
				when 16#1027# => read_data_o <= x"0000";
				when 16#1028# => read_data_o <= x"0000";
				when 16#1029# => read_data_o <= x"0000";
				when 16#102a# => read_data_o <= x"0000";
				when 16#102b# => read_data_o <= x"0000";
				when 16#102c# => read_data_o <= x"0000";
				when 16#102d# => read_data_o <= x"0000";
				when 16#102e# => read_data_o <= x"0000";
				when 16#102f# => read_data_o <= x"0000";
				when 16#1030# => read_data_o <= x"0000";
				when 16#1031# => read_data_o <= x"0000";
				when 16#1032# => read_data_o <= x"0000";
				when 16#1033# => read_data_o <= x"0000";
				when 16#1034# => read_data_o <= x"0000";
				when 16#1035# => read_data_o <= x"0000";
				when 16#1036# => read_data_o <= x"0000";
				when 16#1037# => read_data_o <= x"0000";
				when 16#1038# => read_data_o <= x"0000";
				when 16#1039# => read_data_o <= x"0000";
				when 16#103a# => read_data_o <= x"0000";
				when 16#103b# => read_data_o <= x"0000";
				when 16#103c# => read_data_o <= x"0000";
				when 16#103d# => read_data_o <= x"0000";
				when 16#103e# => read_data_o <= x"0000";
				when 16#103f# => read_data_o <= x"0000";
				when 16#1040# => read_data_o <= x"0000";
				when 16#1041# => read_data_o <= x"0000";
				when 16#1042# => read_data_o <= x"0000";
				when 16#1043# => read_data_o <= x"0000";
				when 16#1044# => read_data_o <= x"0000";
				when 16#1045# => read_data_o <= x"0000";
				when 16#1046# => read_data_o <= x"0000";
				when 16#1047# => read_data_o <= x"0000";
				when 16#1048# => read_data_o <= x"0000";
				when 16#1049# => read_data_o <= x"0000";
				when 16#104a# => read_data_o <= x"0000";
				when 16#104b# => read_data_o <= x"0000";
				when 16#104c# => read_data_o <= x"0000";
				when 16#104d# => read_data_o <= x"0000";
				when 16#104e# => read_data_o <= x"0000";
				when 16#104f# => read_data_o <= x"0000";
				when 16#1050# => read_data_o <= x"0000";
				when 16#1051# => read_data_o <= x"0000";
				when 16#1052# => read_data_o <= x"0000";
				when 16#1053# => read_data_o <= x"0000";
				when 16#1054# => read_data_o <= x"0000";
				when 16#1055# => read_data_o <= x"0000";
				when 16#1056# => read_data_o <= x"0000";
				when 16#1057# => read_data_o <= x"0000";
				when 16#1058# => read_data_o <= x"0000";
				when 16#1059# => read_data_o <= x"0000";
				when 16#105a# => read_data_o <= x"0000";
				when 16#105b# => read_data_o <= x"0000";
				when 16#105c# => read_data_o <= x"0000";
				when 16#105d# => read_data_o <= x"0000";
				when 16#105e# => read_data_o <= x"0000";
				when 16#105f# => read_data_o <= x"0000";
				when 16#1060# => read_data_o <= x"0000";
				when 16#1061# => read_data_o <= x"0000";
				when 16#1062# => read_data_o <= x"0000";
				when 16#1063# => read_data_o <= x"0000";
				when 16#1064# => read_data_o <= x"0000";
				when 16#1065# => read_data_o <= x"0000";
				when 16#1066# => read_data_o <= x"0000";
				when 16#1067# => read_data_o <= x"0000";
				when 16#1068# => read_data_o <= x"0000";
				when 16#1069# => read_data_o <= x"0000";
				when 16#106a# => read_data_o <= x"0000";
				when 16#106b# => read_data_o <= x"0000";
				when 16#106c# => read_data_o <= x"0000";
				when 16#106d# => read_data_o <= x"0000";
				when 16#106e# => read_data_o <= x"0000";
				when 16#106f# => read_data_o <= x"0000";
				when 16#1070# => read_data_o <= x"0000";
				when 16#1071# => read_data_o <= x"0000";
				when 16#1072# => read_data_o <= x"0000";
				when 16#1073# => read_data_o <= x"0000";
				when 16#1074# => read_data_o <= x"0000";
				when 16#1075# => read_data_o <= x"0000";
				when 16#1076# => read_data_o <= x"0000";
				when 16#1077# => read_data_o <= x"0000";
				when 16#1078# => read_data_o <= x"0000";
				when 16#1079# => read_data_o <= x"0000";
				when 16#107a# => read_data_o <= x"0000";
				when 16#107b# => read_data_o <= x"0000";
				when 16#107c# => read_data_o <= x"0000";
				when 16#107d# => read_data_o <= x"0000";
				when 16#107e# => read_data_o <= x"0000";
				when 16#107f# => read_data_o <= x"0000";
				when 16#1080# => read_data_o <= x"0000";
				when 16#1081# => read_data_o <= x"0000";
				when 16#1082# => read_data_o <= x"0000";
				when 16#1083# => read_data_o <= x"0000";
				when 16#1084# => read_data_o <= x"0000";
				when 16#1085# => read_data_o <= x"0000";
				when 16#1086# => read_data_o <= x"0000";
				when 16#1087# => read_data_o <= x"0000";
				when 16#1088# => read_data_o <= x"0000";
				when 16#1089# => read_data_o <= x"0000";
				when 16#108a# => read_data_o <= x"0000";
				when 16#108b# => read_data_o <= x"0000";
				when 16#108c# => read_data_o <= x"0000";
				when 16#108d# => read_data_o <= x"0000";
				when 16#108e# => read_data_o <= x"0000";
				when 16#108f# => read_data_o <= x"0000";
				when 16#1090# => read_data_o <= x"0000";
				when 16#1091# => read_data_o <= x"0000";
				when 16#1092# => read_data_o <= x"0000";
				when 16#1093# => read_data_o <= x"0000";
				when 16#1094# => read_data_o <= x"0000";
				when 16#1095# => read_data_o <= x"0000";
				when 16#1096# => read_data_o <= x"0000";
				when 16#1097# => read_data_o <= x"0000";
				when 16#1098# => read_data_o <= x"0000";
				when 16#1099# => read_data_o <= x"0000";
				when 16#109a# => read_data_o <= x"0000";
				when 16#109b# => read_data_o <= x"0000";
				when 16#109c# => read_data_o <= x"0000";
				when 16#109d# => read_data_o <= x"0000";
				when 16#109e# => read_data_o <= x"0000";
				when 16#109f# => read_data_o <= x"0000";
				when 16#10a0# => read_data_o <= x"0000";
				when 16#10a1# => read_data_o <= x"0000";
				when 16#10a2# => read_data_o <= x"0000";
				when 16#10a3# => read_data_o <= x"0000";
				when 16#10a4# => read_data_o <= x"0000";
				when 16#10a5# => read_data_o <= x"0000";
				when 16#10a6# => read_data_o <= x"0000";
				when 16#10a7# => read_data_o <= x"0000";
				when 16#10a8# => read_data_o <= x"0000";
				when 16#10a9# => read_data_o <= x"0000";
				when 16#10aa# => read_data_o <= x"0000";
				when 16#10ab# => read_data_o <= x"0000";
				when 16#10ac# => read_data_o <= x"0000";
				when 16#10ad# => read_data_o <= x"0000";
				when 16#10ae# => read_data_o <= x"0000";
				when 16#10af# => read_data_o <= x"0000";
				when 16#10b0# => read_data_o <= x"0000";
				when 16#10b1# => read_data_o <= x"0000";
				when 16#10b2# => read_data_o <= x"0000";
				when 16#10b3# => read_data_o <= x"0000";
				when 16#10b4# => read_data_o <= x"0000";
				when 16#10b5# => read_data_o <= x"0000";
				when 16#10b6# => read_data_o <= x"0000";
				when 16#10b7# => read_data_o <= x"0000";
				when 16#10b8# => read_data_o <= x"0000";
				when 16#10b9# => read_data_o <= x"0000";
				when 16#10ba# => read_data_o <= x"0000";
				when 16#10bb# => read_data_o <= x"0000";
				when 16#10bc# => read_data_o <= x"0000";
				when 16#10bd# => read_data_o <= x"0000";
				when 16#10be# => read_data_o <= x"0000";
				when 16#10bf# => read_data_o <= x"0000";
				when 16#10c0# => read_data_o <= x"0000";
				when 16#10c1# => read_data_o <= x"0000";
				when 16#10c2# => read_data_o <= x"0000";
				when 16#10c3# => read_data_o <= x"0000";
				when 16#10c4# => read_data_o <= x"0000";
				when 16#10c5# => read_data_o <= x"0000";
				when 16#10c6# => read_data_o <= x"0000";
				when 16#10c7# => read_data_o <= x"0000";
				when 16#10c8# => read_data_o <= x"0000";
				when 16#10c9# => read_data_o <= x"0000";
				when 16#10ca# => read_data_o <= x"0000";
				when 16#10cb# => read_data_o <= x"0000";
				when 16#10cc# => read_data_o <= x"0000";
				when 16#10cd# => read_data_o <= x"0000";
				when 16#10ce# => read_data_o <= x"0000";
				when 16#10cf# => read_data_o <= x"0000";
				when 16#10d0# => read_data_o <= x"0000";
				when 16#10d1# => read_data_o <= x"0000";
				when 16#10d2# => read_data_o <= x"0000";
				when 16#10d3# => read_data_o <= x"0000";
				when 16#10d4# => read_data_o <= x"0000";
				when 16#10d5# => read_data_o <= x"0000";
				when 16#10d6# => read_data_o <= x"0000";
				when 16#10d7# => read_data_o <= x"0000";
				when 16#10d8# => read_data_o <= x"0000";
				when 16#10d9# => read_data_o <= x"0000";
				when 16#10da# => read_data_o <= x"0000";
				when 16#10db# => read_data_o <= x"0000";
				when 16#10dc# => read_data_o <= x"0000";
				when 16#10dd# => read_data_o <= x"0000";
				when 16#10de# => read_data_o <= x"0000";
				when 16#10df# => read_data_o <= x"0000";
				when 16#10e0# => read_data_o <= x"0000";
				when 16#10e1# => read_data_o <= x"0000";
				when 16#10e2# => read_data_o <= x"0000";
				when 16#10e3# => read_data_o <= x"0000";
				when 16#10e4# => read_data_o <= x"0000";
				when 16#10e5# => read_data_o <= x"0000";
				when 16#10e6# => read_data_o <= x"0000";
				when 16#10e7# => read_data_o <= x"0000";
				when 16#10e8# => read_data_o <= x"0000";
				when 16#10e9# => read_data_o <= x"0000";
				when 16#10ea# => read_data_o <= x"0000";
				when 16#10eb# => read_data_o <= x"0000";
				when 16#10ec# => read_data_o <= x"0000";
				when 16#10ed# => read_data_o <= x"0000";
				when 16#10ee# => read_data_o <= x"0000";
				when 16#10ef# => read_data_o <= x"0000";
				when 16#10f0# => read_data_o <= x"0000";
				when 16#10f1# => read_data_o <= x"0000";
				when 16#10f2# => read_data_o <= x"0000";
				when 16#10f3# => read_data_o <= x"0000";
				when 16#10f4# => read_data_o <= x"0000";
				when 16#10f5# => read_data_o <= x"0000";
				when 16#10f6# => read_data_o <= x"0000";
				when 16#10f7# => read_data_o <= x"0000";
				when 16#10f8# => read_data_o <= x"0000";
				when 16#10f9# => read_data_o <= x"0000";
				when 16#10fa# => read_data_o <= x"0000";
				when 16#10fb# => read_data_o <= x"0000";
				when 16#10fc# => read_data_o <= x"0000";
				when 16#10fd# => read_data_o <= x"0000";
				when 16#10fe# => read_data_o <= x"0000";
				when 16#10ff# => read_data_o <= x"0000";
				when 16#1100# => read_data_o <= x"0000";
				when 16#1101# => read_data_o <= x"0000";
				when 16#1102# => read_data_o <= x"0000";
				when 16#1103# => read_data_o <= x"0000";
				when 16#1104# => read_data_o <= x"0000";
				when 16#1105# => read_data_o <= x"0000";
				when 16#1106# => read_data_o <= x"0000";
				when 16#1107# => read_data_o <= x"0000";
				when 16#1108# => read_data_o <= x"0000";
				when 16#1109# => read_data_o <= x"0000";
				when 16#110a# => read_data_o <= x"0000";
				when 16#110b# => read_data_o <= x"0000";
				when 16#110c# => read_data_o <= x"0000";
				when 16#110d# => read_data_o <= x"0000";
				when 16#110e# => read_data_o <= x"0000";
				when 16#110f# => read_data_o <= x"0000";
				when 16#1110# => read_data_o <= x"0000";
				when 16#1111# => read_data_o <= x"0000";
				when 16#1112# => read_data_o <= x"0000";
				when 16#1113# => read_data_o <= x"0000";
				when 16#1114# => read_data_o <= x"0000";
				when 16#1115# => read_data_o <= x"0000";
				when 16#1116# => read_data_o <= x"0000";
				when 16#1117# => read_data_o <= x"0000";
				when 16#1118# => read_data_o <= x"0000";
				when 16#1119# => read_data_o <= x"0000";
				when 16#111a# => read_data_o <= x"0000";
				when 16#111b# => read_data_o <= x"0000";
				when 16#111c# => read_data_o <= x"0000";
				when 16#111d# => read_data_o <= x"0000";
				when 16#111e# => read_data_o <= x"0000";
				when 16#111f# => read_data_o <= x"0000";
				when 16#1120# => read_data_o <= x"0000";
				when 16#1121# => read_data_o <= x"0000";
				when 16#1122# => read_data_o <= x"0000";
				when 16#1123# => read_data_o <= x"0000";
				when 16#1124# => read_data_o <= x"0000";
				when 16#1125# => read_data_o <= x"0000";
				when 16#1126# => read_data_o <= x"0000";
				when 16#1127# => read_data_o <= x"0000";
				when 16#1128# => read_data_o <= x"0000";
				when 16#1129# => read_data_o <= x"0000";
				when 16#112a# => read_data_o <= x"0000";
				when 16#112b# => read_data_o <= x"0000";
				when 16#112c# => read_data_o <= x"0000";
				when 16#112d# => read_data_o <= x"0000";
				when 16#112e# => read_data_o <= x"0000";
				when 16#112f# => read_data_o <= x"0000";
				when 16#1130# => read_data_o <= x"0000";
				when 16#1131# => read_data_o <= x"0000";
				when 16#1132# => read_data_o <= x"0000";
				when 16#1133# => read_data_o <= x"0000";
				when 16#1134# => read_data_o <= x"0000";
				when 16#1135# => read_data_o <= x"0000";
				when 16#1136# => read_data_o <= x"0000";
				when 16#1137# => read_data_o <= x"0000";
				when 16#1138# => read_data_o <= x"0000";
				when 16#1139# => read_data_o <= x"0000";
				when 16#113a# => read_data_o <= x"0000";
				when 16#113b# => read_data_o <= x"0000";
				when 16#113c# => read_data_o <= x"0000";
				when 16#113d# => read_data_o <= x"0000";
				when 16#113e# => read_data_o <= x"0000";
				when 16#113f# => read_data_o <= x"0000";
				when 16#1140# => read_data_o <= x"0000";
				when 16#1141# => read_data_o <= x"0000";
				when 16#1142# => read_data_o <= x"0000";
				when 16#1143# => read_data_o <= x"0000";
				when 16#1144# => read_data_o <= x"0000";
				when 16#1145# => read_data_o <= x"0000";
				when 16#1146# => read_data_o <= x"0000";
				when 16#1147# => read_data_o <= x"0000";
				when 16#1148# => read_data_o <= x"0000";
				when 16#1149# => read_data_o <= x"0000";
				when 16#114a# => read_data_o <= x"0000";
				when 16#114b# => read_data_o <= x"0000";
				when 16#114c# => read_data_o <= x"0000";
				when 16#114d# => read_data_o <= x"0000";
				when 16#114e# => read_data_o <= x"0000";
				when 16#114f# => read_data_o <= x"0000";
				when 16#1150# => read_data_o <= x"0000";
				when 16#1151# => read_data_o <= x"0000";
				when 16#1152# => read_data_o <= x"0000";
				when 16#1153# => read_data_o <= x"0000";
				when 16#1154# => read_data_o <= x"0000";
				when 16#1155# => read_data_o <= x"0000";
				when 16#1156# => read_data_o <= x"0000";
				when 16#1157# => read_data_o <= x"0000";
				when 16#1158# => read_data_o <= x"0000";
				when 16#1159# => read_data_o <= x"0000";
				when 16#115a# => read_data_o <= x"0000";
				when 16#115b# => read_data_o <= x"0000";
				when 16#115c# => read_data_o <= x"0000";
				when 16#115d# => read_data_o <= x"0000";
				when 16#115e# => read_data_o <= x"0000";
				when 16#115f# => read_data_o <= x"0000";
				when 16#1160# => read_data_o <= x"0000";
				when 16#1161# => read_data_o <= x"0000";
				when 16#1162# => read_data_o <= x"0000";
				when 16#1163# => read_data_o <= x"0000";
				when 16#1164# => read_data_o <= x"0000";
				when 16#1165# => read_data_o <= x"0000";
				when 16#1166# => read_data_o <= x"0000";
				when 16#1167# => read_data_o <= x"0000";
				when 16#1168# => read_data_o <= x"0000";
				when 16#1169# => read_data_o <= x"0000";
				when 16#116a# => read_data_o <= x"0000";
				when 16#116b# => read_data_o <= x"0000";
				when 16#116c# => read_data_o <= x"0000";
				when 16#116d# => read_data_o <= x"0000";
				when 16#116e# => read_data_o <= x"0000";
				when 16#116f# => read_data_o <= x"0000";
				when 16#1170# => read_data_o <= x"0000";
				when 16#1171# => read_data_o <= x"0000";
				when 16#1172# => read_data_o <= x"0000";
				when 16#1173# => read_data_o <= x"0000";
				when 16#1174# => read_data_o <= x"0000";
				when 16#1175# => read_data_o <= x"0000";
				when 16#1176# => read_data_o <= x"0000";
				when 16#1177# => read_data_o <= x"0000";
				when 16#1178# => read_data_o <= x"0000";
				when 16#1179# => read_data_o <= x"0000";
				when 16#117a# => read_data_o <= x"0000";
				when 16#117b# => read_data_o <= x"0000";
				when 16#117c# => read_data_o <= x"0000";
				when 16#117d# => read_data_o <= x"0000";
				when 16#117e# => read_data_o <= x"0000";
				when 16#117f# => read_data_o <= x"0000";
				when 16#1180# => read_data_o <= x"0000";
				when 16#1181# => read_data_o <= x"0000";
				when 16#1182# => read_data_o <= x"0000";
				when 16#1183# => read_data_o <= x"0000";
				when 16#1184# => read_data_o <= x"0000";
				when 16#1185# => read_data_o <= x"0000";
				when 16#1186# => read_data_o <= x"0000";
				when 16#1187# => read_data_o <= x"0000";
				when 16#1188# => read_data_o <= x"0000";
				when 16#1189# => read_data_o <= x"0000";
				when 16#118a# => read_data_o <= x"0000";
				when 16#118b# => read_data_o <= x"0000";
				when 16#118c# => read_data_o <= x"0000";
				when 16#118d# => read_data_o <= x"0000";
				when 16#118e# => read_data_o <= x"0000";
				when 16#118f# => read_data_o <= x"0000";
				when 16#1190# => read_data_o <= x"0000";
				when 16#1191# => read_data_o <= x"0000";
				when 16#1192# => read_data_o <= x"0000";
				when 16#1193# => read_data_o <= x"0000";
				when 16#1194# => read_data_o <= x"0000";
				when 16#1195# => read_data_o <= x"0000";
				when 16#1196# => read_data_o <= x"0000";
				when 16#1197# => read_data_o <= x"0000";
				when 16#1198# => read_data_o <= x"0000";
				when 16#1199# => read_data_o <= x"0000";
				when 16#119a# => read_data_o <= x"0000";
				when 16#119b# => read_data_o <= x"0000";
				when 16#119c# => read_data_o <= x"0000";
				when 16#119d# => read_data_o <= x"0000";
				when 16#119e# => read_data_o <= x"0000";
				when 16#119f# => read_data_o <= x"0000";
				when 16#11a0# => read_data_o <= x"0000";
				when 16#11a1# => read_data_o <= x"0000";
				when 16#11a2# => read_data_o <= x"0000";
				when 16#11a3# => read_data_o <= x"0000";
				when 16#11a4# => read_data_o <= x"0000";
				when 16#11a5# => read_data_o <= x"0000";
				when 16#11a6# => read_data_o <= x"0000";
				when 16#11a7# => read_data_o <= x"0000";
				when 16#11a8# => read_data_o <= x"0000";
				when 16#11a9# => read_data_o <= x"0000";
				when 16#11aa# => read_data_o <= x"0000";
				when 16#11ab# => read_data_o <= x"0000";
				when 16#11ac# => read_data_o <= x"0000";
				when 16#11ad# => read_data_o <= x"0000";
				when 16#11ae# => read_data_o <= x"0000";
				when 16#11af# => read_data_o <= x"0000";
				when 16#11b0# => read_data_o <= x"0000";
				when 16#11b1# => read_data_o <= x"0000";
				when 16#11b2# => read_data_o <= x"0000";
				when 16#11b3# => read_data_o <= x"0000";
				when 16#11b4# => read_data_o <= x"0000";
				when 16#11b5# => read_data_o <= x"0000";
				when 16#11b6# => read_data_o <= x"0000";
				when 16#11b7# => read_data_o <= x"0000";
				when 16#11b8# => read_data_o <= x"0000";
				when 16#11b9# => read_data_o <= x"0000";
				when 16#11ba# => read_data_o <= x"0000";
				when 16#11bb# => read_data_o <= x"0000";
				when 16#11bc# => read_data_o <= x"0000";
				when 16#11bd# => read_data_o <= x"0000";
				when 16#11be# => read_data_o <= x"0000";
				when 16#11bf# => read_data_o <= x"0000";
				when 16#11c0# => read_data_o <= x"0000";
				when 16#11c1# => read_data_o <= x"0000";
				when 16#11c2# => read_data_o <= x"0000";
				when 16#11c3# => read_data_o <= x"0000";
				when 16#11c4# => read_data_o <= x"0000";
				when 16#11c5# => read_data_o <= x"0000";
				when 16#11c6# => read_data_o <= x"0000";
				when 16#11c7# => read_data_o <= x"0000";
				when 16#11c8# => read_data_o <= x"0000";
				when 16#11c9# => read_data_o <= x"0000";
				when 16#11ca# => read_data_o <= x"0000";
				when 16#11cb# => read_data_o <= x"0000";
				when 16#11cc# => read_data_o <= x"0000";
				when 16#11cd# => read_data_o <= x"0000";
				when 16#11ce# => read_data_o <= x"0000";
				when 16#11cf# => read_data_o <= x"0000";
				when 16#11d0# => read_data_o <= x"0000";
				when 16#11d1# => read_data_o <= x"0000";
				when 16#11d2# => read_data_o <= x"0000";
				when 16#11d3# => read_data_o <= x"0000";
				when 16#11d4# => read_data_o <= x"0000";
				when 16#11d5# => read_data_o <= x"0000";
				when 16#11d6# => read_data_o <= x"0000";
				when 16#11d7# => read_data_o <= x"0000";
				when 16#11d8# => read_data_o <= x"0000";
				when 16#11d9# => read_data_o <= x"0000";
				when 16#11da# => read_data_o <= x"0000";
				when 16#11db# => read_data_o <= x"0000";
				when 16#11dc# => read_data_o <= x"0000";
				when 16#11dd# => read_data_o <= x"0000";
				when 16#11de# => read_data_o <= x"0000";
				when 16#11df# => read_data_o <= x"0000";
				when 16#11e0# => read_data_o <= x"0000";
				when 16#11e1# => read_data_o <= x"0000";
				when 16#11e2# => read_data_o <= x"0000";
				when 16#11e3# => read_data_o <= x"0000";
				when 16#11e4# => read_data_o <= x"0000";
				when 16#11e5# => read_data_o <= x"0000";
				when 16#11e6# => read_data_o <= x"0000";
				when 16#11e7# => read_data_o <= x"0000";
				when 16#11e8# => read_data_o <= x"0000";
				when 16#11e9# => read_data_o <= x"0000";
				when 16#11ea# => read_data_o <= x"0000";
				when 16#11eb# => read_data_o <= x"0000";
				when 16#11ec# => read_data_o <= x"0000";
				when 16#11ed# => read_data_o <= x"0000";
				when 16#11ee# => read_data_o <= x"0000";
				when 16#11ef# => read_data_o <= x"0000";
				when 16#11f0# => read_data_o <= x"0000";
				when 16#11f1# => read_data_o <= x"0000";
				when 16#11f2# => read_data_o <= x"0000";
				when 16#11f3# => read_data_o <= x"0000";
				when 16#11f4# => read_data_o <= x"0000";
				when 16#11f5# => read_data_o <= x"0000";
				when 16#11f6# => read_data_o <= x"0000";
				when 16#11f7# => read_data_o <= x"0000";
				when 16#11f8# => read_data_o <= x"0000";
				when 16#11f9# => read_data_o <= x"0000";
				when 16#11fa# => read_data_o <= x"0000";
				when 16#11fb# => read_data_o <= x"0000";
				when 16#11fc# => read_data_o <= x"0000";
				when 16#11fd# => read_data_o <= x"0000";
				when 16#11fe# => read_data_o <= x"0000";
				when 16#11ff# => read_data_o <= x"0000";
				when 16#1200# => read_data_o <= x"0000";
				when 16#1201# => read_data_o <= x"0000";
				when 16#1202# => read_data_o <= x"0000";
				when 16#1203# => read_data_o <= x"0000";
				when 16#1204# => read_data_o <= x"0000";
				when 16#1205# => read_data_o <= x"0000";
				when 16#1206# => read_data_o <= x"0000";
				when 16#1207# => read_data_o <= x"0000";
				when 16#1208# => read_data_o <= x"0000";
				when 16#1209# => read_data_o <= x"0000";
				when 16#120a# => read_data_o <= x"0000";
				when 16#120b# => read_data_o <= x"0000";
				when 16#120c# => read_data_o <= x"0000";
				when 16#120d# => read_data_o <= x"0000";
				when 16#120e# => read_data_o <= x"0000";
				when 16#120f# => read_data_o <= x"0000";
				when 16#1210# => read_data_o <= x"0000";
				when 16#1211# => read_data_o <= x"0000";
				when 16#1212# => read_data_o <= x"0000";
				when 16#1213# => read_data_o <= x"0000";
				when 16#1214# => read_data_o <= x"0000";
				when 16#1215# => read_data_o <= x"0000";
				when 16#1216# => read_data_o <= x"0000";
				when 16#1217# => read_data_o <= x"0000";
				when 16#1218# => read_data_o <= x"0000";
				when 16#1219# => read_data_o <= x"0000";
				when 16#121a# => read_data_o <= x"0000";
				when 16#121b# => read_data_o <= x"0000";
				when 16#121c# => read_data_o <= x"0000";
				when 16#121d# => read_data_o <= x"0000";
				when 16#121e# => read_data_o <= x"0000";
				when 16#121f# => read_data_o <= x"0000";
				when 16#1220# => read_data_o <= x"0000";
				when 16#1221# => read_data_o <= x"0000";
				when 16#1222# => read_data_o <= x"0000";
				when 16#1223# => read_data_o <= x"0000";
				when 16#1224# => read_data_o <= x"0000";
				when 16#1225# => read_data_o <= x"0000";
				when 16#1226# => read_data_o <= x"0000";
				when 16#1227# => read_data_o <= x"0000";
				when 16#1228# => read_data_o <= x"0000";
				when 16#1229# => read_data_o <= x"0000";
				when 16#122a# => read_data_o <= x"0000";
				when 16#122b# => read_data_o <= x"0000";
				when 16#122c# => read_data_o <= x"0000";
				when 16#122d# => read_data_o <= x"0000";
				when 16#122e# => read_data_o <= x"0000";
				when 16#122f# => read_data_o <= x"0000";
				when 16#1230# => read_data_o <= x"0000";
				when 16#1231# => read_data_o <= x"0000";
				when 16#1232# => read_data_o <= x"0000";
				when 16#1233# => read_data_o <= x"0000";
				when 16#1234# => read_data_o <= x"0000";
				when 16#1235# => read_data_o <= x"0000";
				when 16#1236# => read_data_o <= x"0000";
				when 16#1237# => read_data_o <= x"0000";
				when 16#1238# => read_data_o <= x"0000";
				when 16#1239# => read_data_o <= x"0000";
				when 16#123a# => read_data_o <= x"0000";
				when 16#123b# => read_data_o <= x"0000";
				when 16#123c# => read_data_o <= x"0000";
				when 16#123d# => read_data_o <= x"0000";
				when 16#123e# => read_data_o <= x"0000";
				when 16#123f# => read_data_o <= x"0000";
				when 16#1240# => read_data_o <= x"0000";
				when 16#1241# => read_data_o <= x"0000";
				when 16#1242# => read_data_o <= x"0000";
				when 16#1243# => read_data_o <= x"0000";
				when 16#1244# => read_data_o <= x"0000";
				when 16#1245# => read_data_o <= x"0000";
				when 16#1246# => read_data_o <= x"0000";
				when 16#1247# => read_data_o <= x"0000";
				when 16#1248# => read_data_o <= x"0000";
				when 16#1249# => read_data_o <= x"0000";
				when 16#124a# => read_data_o <= x"0000";
				when 16#124b# => read_data_o <= x"0000";
				when 16#124c# => read_data_o <= x"0000";
				when 16#124d# => read_data_o <= x"0000";
				when 16#124e# => read_data_o <= x"0000";
				when 16#124f# => read_data_o <= x"0000";
				when 16#1250# => read_data_o <= x"0000";
				when 16#1251# => read_data_o <= x"0000";
				when 16#1252# => read_data_o <= x"0000";
				when 16#1253# => read_data_o <= x"0000";
				when 16#1254# => read_data_o <= x"0000";
				when 16#1255# => read_data_o <= x"0000";
				when 16#1256# => read_data_o <= x"0000";
				when 16#1257# => read_data_o <= x"0000";
				when 16#1258# => read_data_o <= x"0000";
				when 16#1259# => read_data_o <= x"0000";
				when 16#125a# => read_data_o <= x"0000";
				when 16#125b# => read_data_o <= x"0000";
				when 16#125c# => read_data_o <= x"0000";
				when 16#125d# => read_data_o <= x"0000";
				when 16#125e# => read_data_o <= x"0000";
				when 16#125f# => read_data_o <= x"0000";
				when 16#1260# => read_data_o <= x"0000";
				when 16#1261# => read_data_o <= x"0000";
				when 16#1262# => read_data_o <= x"0000";
				when 16#1263# => read_data_o <= x"0000";
				when 16#1264# => read_data_o <= x"0000";
				when 16#1265# => read_data_o <= x"0000";
				when 16#1266# => read_data_o <= x"0000";
				when 16#1267# => read_data_o <= x"0000";
				when 16#1268# => read_data_o <= x"0000";
				when 16#1269# => read_data_o <= x"0000";
				when 16#126a# => read_data_o <= x"0000";
				when 16#126b# => read_data_o <= x"0000";
				when 16#126c# => read_data_o <= x"0000";
				when 16#126d# => read_data_o <= x"0000";
				when 16#126e# => read_data_o <= x"0000";
				when 16#126f# => read_data_o <= x"0000";
				when 16#1270# => read_data_o <= x"0000";
				when 16#1271# => read_data_o <= x"0000";
				when 16#1272# => read_data_o <= x"0000";
				when 16#1273# => read_data_o <= x"0000";
				when 16#1274# => read_data_o <= x"0000";
				when 16#1275# => read_data_o <= x"0000";
				when 16#1276# => read_data_o <= x"0000";
				when 16#1277# => read_data_o <= x"0000";
				when 16#1278# => read_data_o <= x"0000";
				when 16#1279# => read_data_o <= x"0000";
				when 16#127a# => read_data_o <= x"0000";
				when 16#127b# => read_data_o <= x"0000";
				when 16#127c# => read_data_o <= x"0000";
				when 16#127d# => read_data_o <= x"0000";
				when 16#127e# => read_data_o <= x"0000";
				when 16#127f# => read_data_o <= x"0000";
				when 16#1280# => read_data_o <= x"0000";
				when 16#1281# => read_data_o <= x"0000";
				when 16#1282# => read_data_o <= x"0000";
				when 16#1283# => read_data_o <= x"0000";
				when 16#1284# => read_data_o <= x"0000";
				when 16#1285# => read_data_o <= x"0000";
				when 16#1286# => read_data_o <= x"0000";
				when 16#1287# => read_data_o <= x"0000";
				when 16#1288# => read_data_o <= x"0000";
				when 16#1289# => read_data_o <= x"0000";
				when 16#128a# => read_data_o <= x"0000";
				when 16#128b# => read_data_o <= x"0000";
				when 16#128c# => read_data_o <= x"0000";
				when 16#128d# => read_data_o <= x"0000";
				when 16#128e# => read_data_o <= x"0000";
				when 16#128f# => read_data_o <= x"0000";
				when 16#1290# => read_data_o <= x"0000";
				when 16#1291# => read_data_o <= x"0000";
				when 16#1292# => read_data_o <= x"0000";
				when 16#1293# => read_data_o <= x"0000";
				when 16#1294# => read_data_o <= x"0000";
				when 16#1295# => read_data_o <= x"0000";
				when 16#1296# => read_data_o <= x"0000";
				when 16#1297# => read_data_o <= x"0000";
				when 16#1298# => read_data_o <= x"0000";
				when 16#1299# => read_data_o <= x"0000";
				when 16#129a# => read_data_o <= x"0000";
				when 16#129b# => read_data_o <= x"0000";
				when 16#129c# => read_data_o <= x"0000";
				when 16#129d# => read_data_o <= x"0000";
				when 16#129e# => read_data_o <= x"0000";
				when 16#129f# => read_data_o <= x"0000";
				when 16#12a0# => read_data_o <= x"0000";
				when 16#12a1# => read_data_o <= x"0000";
				when 16#12a2# => read_data_o <= x"0000";
				when 16#12a3# => read_data_o <= x"0000";
				when 16#12a4# => read_data_o <= x"0000";
				when 16#12a5# => read_data_o <= x"0000";
				when 16#12a6# => read_data_o <= x"0000";
				when 16#12a7# => read_data_o <= x"0000";
				when 16#12a8# => read_data_o <= x"0000";
				when 16#12a9# => read_data_o <= x"0000";
				when 16#12aa# => read_data_o <= x"0000";
				when 16#12ab# => read_data_o <= x"0000";
				when 16#12ac# => read_data_o <= x"0000";
				when 16#12ad# => read_data_o <= x"0000";
				when 16#12ae# => read_data_o <= x"0000";
				when 16#12af# => read_data_o <= x"0000";
				when 16#12b0# => read_data_o <= x"0000";
				when 16#12b1# => read_data_o <= x"0000";
				when 16#12b2# => read_data_o <= x"0000";
				when 16#12b3# => read_data_o <= x"0000";
				when 16#12b4# => read_data_o <= x"0000";
				when 16#12b5# => read_data_o <= x"0000";
				when 16#12b6# => read_data_o <= x"0000";
				when 16#12b7# => read_data_o <= x"0000";
				when 16#12b8# => read_data_o <= x"0000";
				when 16#12b9# => read_data_o <= x"0000";
				when 16#12ba# => read_data_o <= x"0000";
				when 16#12bb# => read_data_o <= x"0000";
				when 16#12bc# => read_data_o <= x"0000";
				when 16#12bd# => read_data_o <= x"0000";
				when 16#12be# => read_data_o <= x"0000";
				when 16#12bf# => read_data_o <= x"0000";
				when 16#12c0# => read_data_o <= x"0000";
				when 16#12c1# => read_data_o <= x"0000";
				when 16#12c2# => read_data_o <= x"0000";
				when 16#12c3# => read_data_o <= x"0000";
				when 16#12c4# => read_data_o <= x"0000";
				when 16#12c5# => read_data_o <= x"0000";
				when 16#12c6# => read_data_o <= x"0000";
				when 16#12c7# => read_data_o <= x"0000";
				when 16#12c8# => read_data_o <= x"0000";
				when 16#12c9# => read_data_o <= x"0000";
				when 16#12ca# => read_data_o <= x"0000";
				when 16#12cb# => read_data_o <= x"0000";
				when 16#12cc# => read_data_o <= x"0000";
				when 16#12cd# => read_data_o <= x"0000";
				when 16#12ce# => read_data_o <= x"0000";
				when 16#12cf# => read_data_o <= x"0000";
				when 16#12d0# => read_data_o <= x"0000";
				when 16#12d1# => read_data_o <= x"0000";
				when 16#12d2# => read_data_o <= x"0000";
				when 16#12d3# => read_data_o <= x"0000";
				when 16#12d4# => read_data_o <= x"0000";
				when 16#12d5# => read_data_o <= x"0000";
				when 16#12d6# => read_data_o <= x"0000";
				when 16#12d7# => read_data_o <= x"0000";
				when 16#12d8# => read_data_o <= x"0000";
				when 16#12d9# => read_data_o <= x"0000";
				when 16#12da# => read_data_o <= x"0000";
				when 16#12db# => read_data_o <= x"0000";
				when 16#12dc# => read_data_o <= x"0000";
				when 16#12dd# => read_data_o <= x"0000";
				when 16#12de# => read_data_o <= x"0000";
				when 16#12df# => read_data_o <= x"0000";
				when 16#12e0# => read_data_o <= x"0000";
				when 16#12e1# => read_data_o <= x"0000";
				when 16#12e2# => read_data_o <= x"0000";
				when 16#12e3# => read_data_o <= x"0000";
				when 16#12e4# => read_data_o <= x"0000";
				when 16#12e5# => read_data_o <= x"0000";
				when 16#12e6# => read_data_o <= x"0000";
				when 16#12e7# => read_data_o <= x"0000";
				when 16#12e8# => read_data_o <= x"0000";
				when 16#12e9# => read_data_o <= x"0000";
				when 16#12ea# => read_data_o <= x"0000";
				when 16#12eb# => read_data_o <= x"0000";
				when 16#12ec# => read_data_o <= x"0000";
				when 16#12ed# => read_data_o <= x"0000";
				when 16#12ee# => read_data_o <= x"0000";
				when 16#12ef# => read_data_o <= x"0000";
				when 16#12f0# => read_data_o <= x"0000";
				when 16#12f1# => read_data_o <= x"0000";
				when 16#12f2# => read_data_o <= x"0000";
				when 16#12f3# => read_data_o <= x"0000";
				when 16#12f4# => read_data_o <= x"0000";
				when 16#12f5# => read_data_o <= x"0000";
				when 16#12f6# => read_data_o <= x"0000";
				when 16#12f7# => read_data_o <= x"0000";
				when 16#12f8# => read_data_o <= x"0000";
				when 16#12f9# => read_data_o <= x"0000";
				when 16#12fa# => read_data_o <= x"0000";
				when 16#12fb# => read_data_o <= x"0000";
				when 16#12fc# => read_data_o <= x"0000";
				when 16#12fd# => read_data_o <= x"0000";
				when 16#12fe# => read_data_o <= x"0000";
				when 16#12ff# => read_data_o <= x"0000";
				when 16#1300# => read_data_o <= x"0000";
				when 16#1301# => read_data_o <= x"0000";
				when 16#1302# => read_data_o <= x"0000";
				when 16#1303# => read_data_o <= x"0000";
				when 16#1304# => read_data_o <= x"0000";
				when 16#1305# => read_data_o <= x"0000";
				when 16#1306# => read_data_o <= x"0000";
				when 16#1307# => read_data_o <= x"0000";
				when 16#1308# => read_data_o <= x"0000";
				when 16#1309# => read_data_o <= x"0000";
				when 16#130a# => read_data_o <= x"0000";
				when 16#130b# => read_data_o <= x"0000";
				when 16#130c# => read_data_o <= x"0000";
				when 16#130d# => read_data_o <= x"0000";
				when 16#130e# => read_data_o <= x"0000";
				when 16#130f# => read_data_o <= x"0000";
				when 16#1310# => read_data_o <= x"0000";
				when 16#1311# => read_data_o <= x"0000";
				when 16#1312# => read_data_o <= x"0000";
				when 16#1313# => read_data_o <= x"0000";
				when 16#1314# => read_data_o <= x"0000";
				when 16#1315# => read_data_o <= x"0000";
				when 16#1316# => read_data_o <= x"0000";
				when 16#1317# => read_data_o <= x"0000";
				when 16#1318# => read_data_o <= x"0000";
				when 16#1319# => read_data_o <= x"0000";
				when 16#131a# => read_data_o <= x"0000";
				when 16#131b# => read_data_o <= x"0000";
				when 16#131c# => read_data_o <= x"0000";
				when 16#131d# => read_data_o <= x"0000";
				when 16#131e# => read_data_o <= x"0000";
				when 16#131f# => read_data_o <= x"0000";
				when 16#1320# => read_data_o <= x"0000";
				when 16#1321# => read_data_o <= x"0000";
				when 16#1322# => read_data_o <= x"0000";
				when 16#1323# => read_data_o <= x"0000";
				when 16#1324# => read_data_o <= x"0000";
				when 16#1325# => read_data_o <= x"0000";
				when 16#1326# => read_data_o <= x"0000";
				when 16#1327# => read_data_o <= x"0000";
				when 16#1328# => read_data_o <= x"0000";
				when 16#1329# => read_data_o <= x"0000";
				when 16#132a# => read_data_o <= x"0000";
				when 16#132b# => read_data_o <= x"0000";
				when 16#132c# => read_data_o <= x"0000";
				when 16#132d# => read_data_o <= x"0000";
				when 16#132e# => read_data_o <= x"0000";
				when 16#132f# => read_data_o <= x"0000";
				when 16#1330# => read_data_o <= x"0000";
				when 16#1331# => read_data_o <= x"0000";
				when 16#1332# => read_data_o <= x"0000";
				when 16#1333# => read_data_o <= x"0000";
				when 16#1334# => read_data_o <= x"0000";
				when 16#1335# => read_data_o <= x"0000";
				when 16#1336# => read_data_o <= x"0000";
				when 16#1337# => read_data_o <= x"0000";
				when 16#1338# => read_data_o <= x"0000";
				when 16#1339# => read_data_o <= x"0000";
				when 16#133a# => read_data_o <= x"0000";
				when 16#133b# => read_data_o <= x"0000";
				when 16#133c# => read_data_o <= x"0000";
				when 16#133d# => read_data_o <= x"0000";
				when 16#133e# => read_data_o <= x"0000";
				when 16#133f# => read_data_o <= x"0000";
				when 16#1340# => read_data_o <= x"0000";
				when 16#1341# => read_data_o <= x"0000";
				when 16#1342# => read_data_o <= x"0000";
				when 16#1343# => read_data_o <= x"0000";
				when 16#1344# => read_data_o <= x"0000";
				when 16#1345# => read_data_o <= x"0000";
				when 16#1346# => read_data_o <= x"0000";
				when 16#1347# => read_data_o <= x"0000";
				when 16#1348# => read_data_o <= x"0000";
				when 16#1349# => read_data_o <= x"0000";
				when 16#134a# => read_data_o <= x"0000";
				when 16#134b# => read_data_o <= x"0000";
				when 16#134c# => read_data_o <= x"0000";
				when 16#134d# => read_data_o <= x"0000";
				when 16#134e# => read_data_o <= x"0000";
				when 16#134f# => read_data_o <= x"0000";
				when 16#1350# => read_data_o <= x"0000";
				when 16#1351# => read_data_o <= x"0000";
				when 16#1352# => read_data_o <= x"0000";
				when 16#1353# => read_data_o <= x"0000";
				when 16#1354# => read_data_o <= x"0000";
				when 16#1355# => read_data_o <= x"0000";
				when 16#1356# => read_data_o <= x"0000";
				when 16#1357# => read_data_o <= x"0000";
				when 16#1358# => read_data_o <= x"0000";
				when 16#1359# => read_data_o <= x"0000";
				when 16#135a# => read_data_o <= x"0000";
				when 16#135b# => read_data_o <= x"0000";
				when 16#135c# => read_data_o <= x"0000";
				when 16#135d# => read_data_o <= x"0000";
				when 16#135e# => read_data_o <= x"0000";
				when 16#135f# => read_data_o <= x"0000";
				when 16#1360# => read_data_o <= x"0000";
				when 16#1361# => read_data_o <= x"0000";
				when 16#1362# => read_data_o <= x"0000";
				when 16#1363# => read_data_o <= x"0000";
				when 16#1364# => read_data_o <= x"0000";
				when 16#1365# => read_data_o <= x"0000";
				when 16#1366# => read_data_o <= x"0000";
				when 16#1367# => read_data_o <= x"0000";
				when 16#1368# => read_data_o <= x"0000";
				when 16#1369# => read_data_o <= x"0000";
				when 16#136a# => read_data_o <= x"0000";
				when 16#136b# => read_data_o <= x"0000";
				when 16#136c# => read_data_o <= x"0000";
				when 16#136d# => read_data_o <= x"0000";
				when 16#136e# => read_data_o <= x"0000";
				when 16#136f# => read_data_o <= x"0000";
				when 16#1370# => read_data_o <= x"0000";
				when 16#1371# => read_data_o <= x"0000";
				when 16#1372# => read_data_o <= x"0000";
				when 16#1373# => read_data_o <= x"0000";
				when 16#1374# => read_data_o <= x"0000";
				when 16#1375# => read_data_o <= x"0000";
				when 16#1376# => read_data_o <= x"0000";
				when 16#1377# => read_data_o <= x"0000";
				when 16#1378# => read_data_o <= x"0000";
				when 16#1379# => read_data_o <= x"0000";
				when 16#137a# => read_data_o <= x"0000";
				when 16#137b# => read_data_o <= x"0000";
				when 16#137c# => read_data_o <= x"0000";
				when 16#137d# => read_data_o <= x"0000";
				when 16#137e# => read_data_o <= x"0000";
				when 16#137f# => read_data_o <= x"0000";
				when 16#1380# => read_data_o <= x"0000";
				when 16#1381# => read_data_o <= x"0000";
				when 16#1382# => read_data_o <= x"0000";
				when 16#1383# => read_data_o <= x"0000";
				when 16#1384# => read_data_o <= x"0000";
				when 16#1385# => read_data_o <= x"0000";
				when 16#1386# => read_data_o <= x"0000";
				when 16#1387# => read_data_o <= x"0000";
				when 16#1388# => read_data_o <= x"0000";
				when 16#1389# => read_data_o <= x"0000";
				when 16#138a# => read_data_o <= x"0000";
				when 16#138b# => read_data_o <= x"0000";
				when 16#138c# => read_data_o <= x"0000";
				when 16#138d# => read_data_o <= x"0000";
				when 16#138e# => read_data_o <= x"0000";
				when 16#138f# => read_data_o <= x"0000";
				when 16#1390# => read_data_o <= x"0000";
				when 16#1391# => read_data_o <= x"0000";
				when 16#1392# => read_data_o <= x"0000";
				when 16#1393# => read_data_o <= x"0000";
				when 16#1394# => read_data_o <= x"0000";
				when 16#1395# => read_data_o <= x"0000";
				when 16#1396# => read_data_o <= x"0000";
				when 16#1397# => read_data_o <= x"0000";
				when 16#1398# => read_data_o <= x"0000";
				when 16#1399# => read_data_o <= x"0000";
				when 16#139a# => read_data_o <= x"0000";
				when 16#139b# => read_data_o <= x"0000";
				when 16#139c# => read_data_o <= x"0000";
				when 16#139d# => read_data_o <= x"0000";
				when 16#139e# => read_data_o <= x"0000";
				when 16#139f# => read_data_o <= x"0000";
				when 16#13a0# => read_data_o <= x"0000";
				when 16#13a1# => read_data_o <= x"0000";
				when 16#13a2# => read_data_o <= x"0000";
				when 16#13a3# => read_data_o <= x"0000";
				when 16#13a4# => read_data_o <= x"0000";
				when 16#13a5# => read_data_o <= x"0000";
				when 16#13a6# => read_data_o <= x"0000";
				when 16#13a7# => read_data_o <= x"0000";
				when 16#13a8# => read_data_o <= x"0000";
				when 16#13a9# => read_data_o <= x"0000";
				when 16#13aa# => read_data_o <= x"0000";
				when 16#13ab# => read_data_o <= x"0000";
				when 16#13ac# => read_data_o <= x"0000";
				when 16#13ad# => read_data_o <= x"0000";
				when 16#13ae# => read_data_o <= x"0000";
				when 16#13af# => read_data_o <= x"0000";
				when 16#13b0# => read_data_o <= x"0000";
				when 16#13b1# => read_data_o <= x"0000";
				when 16#13b2# => read_data_o <= x"0000";
				when 16#13b3# => read_data_o <= x"0000";
				when 16#13b4# => read_data_o <= x"0000";
				when 16#13b5# => read_data_o <= x"0000";
				when 16#13b6# => read_data_o <= x"0000";
				when 16#13b7# => read_data_o <= x"0000";
				when 16#13b8# => read_data_o <= x"0000";
				when 16#13b9# => read_data_o <= x"0000";
				when 16#13ba# => read_data_o <= x"0000";
				when 16#13bb# => read_data_o <= x"0000";
				when 16#13bc# => read_data_o <= x"0000";
				when 16#13bd# => read_data_o <= x"0000";
				when 16#13be# => read_data_o <= x"0000";
				when 16#13bf# => read_data_o <= x"0000";
				when 16#13c0# => read_data_o <= x"0000";
				when 16#13c1# => read_data_o <= x"0000";
				when 16#13c2# => read_data_o <= x"0000";
				when 16#13c3# => read_data_o <= x"0000";
				when 16#13c4# => read_data_o <= x"0000";
				when 16#13c5# => read_data_o <= x"0000";
				when 16#13c6# => read_data_o <= x"0000";
				when 16#13c7# => read_data_o <= x"0000";
				when 16#13c8# => read_data_o <= x"0000";
				when 16#13c9# => read_data_o <= x"0000";
				when 16#13ca# => read_data_o <= x"0000";
				when 16#13cb# => read_data_o <= x"0000";
				when 16#13cc# => read_data_o <= x"0000";
				when 16#13cd# => read_data_o <= x"0000";
				when 16#13ce# => read_data_o <= x"0000";
				when 16#13cf# => read_data_o <= x"0000";
				when 16#13d0# => read_data_o <= x"0000";
				when 16#13d1# => read_data_o <= x"0000";
				when 16#13d2# => read_data_o <= x"0000";
				when 16#13d3# => read_data_o <= x"0000";
				when 16#13d4# => read_data_o <= x"0000";
				when 16#13d5# => read_data_o <= x"0000";
				when 16#13d6# => read_data_o <= x"0000";
				when 16#13d7# => read_data_o <= x"0000";
				when 16#13d8# => read_data_o <= x"0000";
				when 16#13d9# => read_data_o <= x"0000";
				when 16#13da# => read_data_o <= x"0000";
				when 16#13db# => read_data_o <= x"0000";
				when 16#13dc# => read_data_o <= x"0000";
				when 16#13dd# => read_data_o <= x"0000";
				when 16#13de# => read_data_o <= x"0000";
				when 16#13df# => read_data_o <= x"0000";
				when 16#13e0# => read_data_o <= x"0000";
				when 16#13e1# => read_data_o <= x"0000";
				when 16#13e2# => read_data_o <= x"0000";
				when 16#13e3# => read_data_o <= x"0000";
				when 16#13e4# => read_data_o <= x"0000";
				when 16#13e5# => read_data_o <= x"0000";
				when 16#13e6# => read_data_o <= x"0000";
				when 16#13e7# => read_data_o <= x"0000";
				when 16#13e8# => read_data_o <= x"0000";
				when 16#13e9# => read_data_o <= x"0000";
				when 16#13ea# => read_data_o <= x"0000";
				when 16#13eb# => read_data_o <= x"0000";
				when 16#13ec# => read_data_o <= x"0000";
				when 16#13ed# => read_data_o <= x"0000";
				when 16#13ee# => read_data_o <= x"0000";
				when 16#13ef# => read_data_o <= x"0000";
				when 16#13f0# => read_data_o <= x"0000";
				when 16#13f1# => read_data_o <= x"0000";
				when 16#13f2# => read_data_o <= x"0000";
				when 16#13f3# => read_data_o <= x"0000";
				when 16#13f4# => read_data_o <= x"0000";
				when 16#13f5# => read_data_o <= x"0000";
				when 16#13f6# => read_data_o <= x"0000";
				when 16#13f7# => read_data_o <= x"0000";
				when 16#13f8# => read_data_o <= x"0000";
				when 16#13f9# => read_data_o <= x"0000";
				when 16#13fa# => read_data_o <= x"0000";
				when 16#13fb# => read_data_o <= x"0000";
				when 16#13fc# => read_data_o <= x"0000";
				when 16#13fd# => read_data_o <= x"0000";
				when 16#13fe# => read_data_o <= x"0000";
				when 16#13ff# => read_data_o <= x"0000";
				when 16#1400# => read_data_o <= x"0000";
				when 16#1401# => read_data_o <= x"0000";
				when 16#1402# => read_data_o <= x"0000";
				when 16#1403# => read_data_o <= x"0000";
				when 16#1404# => read_data_o <= x"0000";
				when 16#1405# => read_data_o <= x"0000";
				when 16#1406# => read_data_o <= x"0000";
				when 16#1407# => read_data_o <= x"0000";
				when 16#1408# => read_data_o <= x"0000";
				when 16#1409# => read_data_o <= x"0000";
				when 16#140a# => read_data_o <= x"0000";
				when 16#140b# => read_data_o <= x"0000";
				when 16#140c# => read_data_o <= x"0000";
				when 16#140d# => read_data_o <= x"0000";
				when 16#140e# => read_data_o <= x"0000";
				when 16#140f# => read_data_o <= x"0000";
				when 16#1410# => read_data_o <= x"0000";
				when 16#1411# => read_data_o <= x"0000";
				when 16#1412# => read_data_o <= x"0000";
				when 16#1413# => read_data_o <= x"0000";
				when 16#1414# => read_data_o <= x"0000";
				when 16#1415# => read_data_o <= x"0000";
				when 16#1416# => read_data_o <= x"0000";
				when 16#1417# => read_data_o <= x"0000";
				when 16#1418# => read_data_o <= x"0000";
				when 16#1419# => read_data_o <= x"0000";
				when 16#141a# => read_data_o <= x"0000";
				when 16#141b# => read_data_o <= x"0000";
				when 16#141c# => read_data_o <= x"0000";
				when 16#141d# => read_data_o <= x"0000";
				when 16#141e# => read_data_o <= x"0000";
				when 16#141f# => read_data_o <= x"0000";
				when 16#1420# => read_data_o <= x"0000";
				when 16#1421# => read_data_o <= x"0000";
				when 16#1422# => read_data_o <= x"0000";
				when 16#1423# => read_data_o <= x"0000";
				when 16#1424# => read_data_o <= x"0000";
				when 16#1425# => read_data_o <= x"0000";
				when 16#1426# => read_data_o <= x"0000";
				when 16#1427# => read_data_o <= x"0000";
				when 16#1428# => read_data_o <= x"0000";
				when 16#1429# => read_data_o <= x"0000";
				when 16#142a# => read_data_o <= x"0000";
				when 16#142b# => read_data_o <= x"0000";
				when 16#142c# => read_data_o <= x"0000";
				when 16#142d# => read_data_o <= x"0000";
				when 16#142e# => read_data_o <= x"0000";
				when 16#142f# => read_data_o <= x"0000";
				when 16#1430# => read_data_o <= x"0000";
				when 16#1431# => read_data_o <= x"0000";
				when 16#1432# => read_data_o <= x"0000";
				when 16#1433# => read_data_o <= x"0000";
				when 16#1434# => read_data_o <= x"0000";
				when 16#1435# => read_data_o <= x"0000";
				when 16#1436# => read_data_o <= x"0000";
				when 16#1437# => read_data_o <= x"0000";
				when 16#1438# => read_data_o <= x"0000";
				when 16#1439# => read_data_o <= x"0000";
				when 16#143a# => read_data_o <= x"0000";
				when 16#143b# => read_data_o <= x"0000";
				when 16#143c# => read_data_o <= x"0000";
				when 16#143d# => read_data_o <= x"0000";
				when 16#143e# => read_data_o <= x"0000";
				when 16#143f# => read_data_o <= x"0000";
				when 16#1440# => read_data_o <= x"0000";
				when 16#1441# => read_data_o <= x"0000";
				when 16#1442# => read_data_o <= x"0000";
				when 16#1443# => read_data_o <= x"0000";
				when 16#1444# => read_data_o <= x"0000";
				when 16#1445# => read_data_o <= x"0000";
				when 16#1446# => read_data_o <= x"0000";
				when 16#1447# => read_data_o <= x"0000";
				when 16#1448# => read_data_o <= x"0000";
				when 16#1449# => read_data_o <= x"0000";
				when 16#144a# => read_data_o <= x"0000";
				when 16#144b# => read_data_o <= x"0000";
				when 16#144c# => read_data_o <= x"0000";
				when 16#144d# => read_data_o <= x"0000";
				when 16#144e# => read_data_o <= x"0000";
				when 16#144f# => read_data_o <= x"0000";
				when 16#1450# => read_data_o <= x"0000";
				when 16#1451# => read_data_o <= x"0000";
				when 16#1452# => read_data_o <= x"0000";
				when 16#1453# => read_data_o <= x"0000";
				when 16#1454# => read_data_o <= x"0000";
				when 16#1455# => read_data_o <= x"0000";
				when 16#1456# => read_data_o <= x"0000";
				when 16#1457# => read_data_o <= x"0000";
				when 16#1458# => read_data_o <= x"0000";
				when 16#1459# => read_data_o <= x"0000";
				when 16#145a# => read_data_o <= x"0000";
				when 16#145b# => read_data_o <= x"0000";
				when 16#145c# => read_data_o <= x"0000";
				when 16#145d# => read_data_o <= x"0000";
				when 16#145e# => read_data_o <= x"0000";
				when 16#145f# => read_data_o <= x"0000";
				when 16#1460# => read_data_o <= x"0000";
				when 16#1461# => read_data_o <= x"0000";
				when 16#1462# => read_data_o <= x"0000";
				when 16#1463# => read_data_o <= x"0000";
				when 16#1464# => read_data_o <= x"0000";
				when 16#1465# => read_data_o <= x"0000";
				when 16#1466# => read_data_o <= x"0000";
				when 16#1467# => read_data_o <= x"0000";
				when 16#1468# => read_data_o <= x"0000";
				when 16#1469# => read_data_o <= x"0000";
				when 16#146a# => read_data_o <= x"0000";
				when 16#146b# => read_data_o <= x"0000";
				when 16#146c# => read_data_o <= x"0000";
				when 16#146d# => read_data_o <= x"0000";
				when 16#146e# => read_data_o <= x"0000";
				when 16#146f# => read_data_o <= x"0000";
				when 16#1470# => read_data_o <= x"0000";
				when 16#1471# => read_data_o <= x"0000";
				when 16#1472# => read_data_o <= x"0000";
				when 16#1473# => read_data_o <= x"0000";
				when 16#1474# => read_data_o <= x"0000";
				when 16#1475# => read_data_o <= x"0000";
				when 16#1476# => read_data_o <= x"0000";
				when 16#1477# => read_data_o <= x"0000";
				when 16#1478# => read_data_o <= x"0000";
				when 16#1479# => read_data_o <= x"0000";
				when 16#147a# => read_data_o <= x"0000";
				when 16#147b# => read_data_o <= x"0000";
				when 16#147c# => read_data_o <= x"0000";
				when 16#147d# => read_data_o <= x"0000";
				when 16#147e# => read_data_o <= x"0000";
				when 16#147f# => read_data_o <= x"0000";
				when 16#1480# => read_data_o <= x"0000";
				when 16#1481# => read_data_o <= x"0000";
				when 16#1482# => read_data_o <= x"0000";
				when 16#1483# => read_data_o <= x"0000";
				when 16#1484# => read_data_o <= x"0000";
				when 16#1485# => read_data_o <= x"0000";
				when 16#1486# => read_data_o <= x"0000";
				when 16#1487# => read_data_o <= x"0000";
				when 16#1488# => read_data_o <= x"0000";
				when 16#1489# => read_data_o <= x"0000";
				when 16#148a# => read_data_o <= x"0000";
				when 16#148b# => read_data_o <= x"0000";
				when 16#148c# => read_data_o <= x"0000";
				when 16#148d# => read_data_o <= x"0000";
				when 16#148e# => read_data_o <= x"0000";
				when 16#148f# => read_data_o <= x"0000";
				when 16#1490# => read_data_o <= x"0000";
				when 16#1491# => read_data_o <= x"0000";
				when 16#1492# => read_data_o <= x"0000";
				when 16#1493# => read_data_o <= x"0000";
				when 16#1494# => read_data_o <= x"0000";
				when 16#1495# => read_data_o <= x"0000";
				when 16#1496# => read_data_o <= x"0000";
				when 16#1497# => read_data_o <= x"0000";
				when 16#1498# => read_data_o <= x"0000";
				when 16#1499# => read_data_o <= x"0000";
				when 16#149a# => read_data_o <= x"0000";
				when 16#149b# => read_data_o <= x"0000";
				when 16#149c# => read_data_o <= x"0000";
				when 16#149d# => read_data_o <= x"0000";
				when 16#149e# => read_data_o <= x"0000";
				when 16#149f# => read_data_o <= x"0000";
				when 16#14a0# => read_data_o <= x"0000";
				when 16#14a1# => read_data_o <= x"0000";
				when 16#14a2# => read_data_o <= x"0000";
				when 16#14a3# => read_data_o <= x"0000";
				when 16#14a4# => read_data_o <= x"0000";
				when 16#14a5# => read_data_o <= x"0000";
				when 16#14a6# => read_data_o <= x"0000";
				when 16#14a7# => read_data_o <= x"0000";
				when 16#14a8# => read_data_o <= x"0000";
				when 16#14a9# => read_data_o <= x"0000";
				when 16#14aa# => read_data_o <= x"0000";
				when 16#14ab# => read_data_o <= x"0000";
				when 16#14ac# => read_data_o <= x"0000";
				when 16#14ad# => read_data_o <= x"0000";
				when 16#14ae# => read_data_o <= x"0000";
				when 16#14af# => read_data_o <= x"0000";
				when 16#14b0# => read_data_o <= x"0000";
				when 16#14b1# => read_data_o <= x"0000";
				when 16#14b2# => read_data_o <= x"0000";
				when 16#14b3# => read_data_o <= x"0000";
				when 16#14b4# => read_data_o <= x"0000";
				when 16#14b5# => read_data_o <= x"0000";
				when 16#14b6# => read_data_o <= x"0000";
				when 16#14b7# => read_data_o <= x"0000";
				when 16#14b8# => read_data_o <= x"0000";
				when 16#14b9# => read_data_o <= x"0000";
				when 16#14ba# => read_data_o <= x"0000";
				when 16#14bb# => read_data_o <= x"0000";
				when 16#14bc# => read_data_o <= x"0000";
				when 16#14bd# => read_data_o <= x"0000";
				when 16#14be# => read_data_o <= x"0000";
				when 16#14bf# => read_data_o <= x"0000";
				when 16#14c0# => read_data_o <= x"0000";
				when 16#14c1# => read_data_o <= x"0000";
				when 16#14c2# => read_data_o <= x"0000";
				when 16#14c3# => read_data_o <= x"0000";
				when 16#14c4# => read_data_o <= x"0000";
				when 16#14c5# => read_data_o <= x"0000";
				when 16#14c6# => read_data_o <= x"0000";
				when 16#14c7# => read_data_o <= x"0000";
				when 16#14c8# => read_data_o <= x"0000";
				when 16#14c9# => read_data_o <= x"0000";
				when 16#14ca# => read_data_o <= x"0000";
				when 16#14cb# => read_data_o <= x"0000";
				when 16#14cc# => read_data_o <= x"0000";
				when 16#14cd# => read_data_o <= x"0000";
				when 16#14ce# => read_data_o <= x"0000";
				when 16#14cf# => read_data_o <= x"0000";
				when 16#14d0# => read_data_o <= x"0000";
				when 16#14d1# => read_data_o <= x"0000";
				when 16#14d2# => read_data_o <= x"0000";
				when 16#14d3# => read_data_o <= x"0000";
				when 16#14d4# => read_data_o <= x"0000";
				when 16#14d5# => read_data_o <= x"0000";
				when 16#14d6# => read_data_o <= x"0000";
				when 16#14d7# => read_data_o <= x"0000";
				when 16#14d8# => read_data_o <= x"0000";
				when 16#14d9# => read_data_o <= x"0000";
				when 16#14da# => read_data_o <= x"0000";
				when 16#14db# => read_data_o <= x"0000";
				when 16#14dc# => read_data_o <= x"0000";
				when 16#14dd# => read_data_o <= x"0000";
				when 16#14de# => read_data_o <= x"0000";
				when 16#14df# => read_data_o <= x"0000";
				when 16#14e0# => read_data_o <= x"0000";
				when 16#14e1# => read_data_o <= x"0000";
				when 16#14e2# => read_data_o <= x"0000";
				when 16#14e3# => read_data_o <= x"0000";
				when 16#14e4# => read_data_o <= x"0000";
				when 16#14e5# => read_data_o <= x"0000";
				when 16#14e6# => read_data_o <= x"0000";
				when 16#14e7# => read_data_o <= x"0000";
				when 16#14e8# => read_data_o <= x"0000";
				when 16#14e9# => read_data_o <= x"0000";
				when 16#14ea# => read_data_o <= x"0000";
				when 16#14eb# => read_data_o <= x"0000";
				when 16#14ec# => read_data_o <= x"0000";
				when 16#14ed# => read_data_o <= x"0000";
				when 16#14ee# => read_data_o <= x"0000";
				when 16#14ef# => read_data_o <= x"0000";
				when 16#14f0# => read_data_o <= x"0000";
				when 16#14f1# => read_data_o <= x"0000";
				when 16#14f2# => read_data_o <= x"0000";
				when 16#14f3# => read_data_o <= x"0000";
				when 16#14f4# => read_data_o <= x"0000";
				when 16#14f5# => read_data_o <= x"0000";
				when 16#14f6# => read_data_o <= x"0000";
				when 16#14f7# => read_data_o <= x"0000";
				when 16#14f8# => read_data_o <= x"0000";
				when 16#14f9# => read_data_o <= x"0000";
				when 16#14fa# => read_data_o <= x"0000";
				when 16#14fb# => read_data_o <= x"0000";
				when 16#14fc# => read_data_o <= x"0000";
				when 16#14fd# => read_data_o <= x"0000";
				when 16#14fe# => read_data_o <= x"0000";
				when 16#14ff# => read_data_o <= x"0000";
				when 16#1500# => read_data_o <= x"0000";
				when 16#1501# => read_data_o <= x"0000";
				when 16#1502# => read_data_o <= x"0000";
				when 16#1503# => read_data_o <= x"0000";
				when 16#1504# => read_data_o <= x"0000";
				when 16#1505# => read_data_o <= x"0000";
				when 16#1506# => read_data_o <= x"0000";
				when 16#1507# => read_data_o <= x"0000";
				when 16#1508# => read_data_o <= x"0000";
				when 16#1509# => read_data_o <= x"0000";
				when 16#150a# => read_data_o <= x"0000";
				when 16#150b# => read_data_o <= x"0000";
				when 16#150c# => read_data_o <= x"0000";
				when 16#150d# => read_data_o <= x"0000";
				when 16#150e# => read_data_o <= x"0000";
				when 16#150f# => read_data_o <= x"0000";
				when 16#1510# => read_data_o <= x"0000";
				when 16#1511# => read_data_o <= x"0000";
				when 16#1512# => read_data_o <= x"0000";
				when 16#1513# => read_data_o <= x"0000";
				when 16#1514# => read_data_o <= x"0000";
				when 16#1515# => read_data_o <= x"0000";
				when 16#1516# => read_data_o <= x"0000";
				when 16#1517# => read_data_o <= x"0000";
				when 16#1518# => read_data_o <= x"0000";
				when 16#1519# => read_data_o <= x"0000";
				when 16#151a# => read_data_o <= x"0000";
				when 16#151b# => read_data_o <= x"0000";
				when 16#151c# => read_data_o <= x"0000";
				when 16#151d# => read_data_o <= x"0000";
				when 16#151e# => read_data_o <= x"0000";
				when 16#151f# => read_data_o <= x"0000";
				when 16#1520# => read_data_o <= x"0000";
				when 16#1521# => read_data_o <= x"0000";
				when 16#1522# => read_data_o <= x"0000";
				when 16#1523# => read_data_o <= x"0000";
				when 16#1524# => read_data_o <= x"0000";
				when 16#1525# => read_data_o <= x"0000";
				when 16#1526# => read_data_o <= x"0000";
				when 16#1527# => read_data_o <= x"0000";
				when 16#1528# => read_data_o <= x"0000";
				when 16#1529# => read_data_o <= x"0000";
				when 16#152a# => read_data_o <= x"0000";
				when 16#152b# => read_data_o <= x"0000";
				when 16#152c# => read_data_o <= x"0000";
				when 16#152d# => read_data_o <= x"0000";
				when 16#152e# => read_data_o <= x"0000";
				when 16#152f# => read_data_o <= x"0000";
				when 16#1530# => read_data_o <= x"0000";
				when 16#1531# => read_data_o <= x"0000";
				when 16#1532# => read_data_o <= x"0000";
				when 16#1533# => read_data_o <= x"0000";
				when 16#1534# => read_data_o <= x"0000";
				when 16#1535# => read_data_o <= x"0000";
				when 16#1536# => read_data_o <= x"0000";
				when 16#1537# => read_data_o <= x"0000";
				when 16#1538# => read_data_o <= x"0000";
				when 16#1539# => read_data_o <= x"0000";
				when 16#153a# => read_data_o <= x"0000";
				when 16#153b# => read_data_o <= x"0000";
				when 16#153c# => read_data_o <= x"0000";
				when 16#153d# => read_data_o <= x"0000";
				when 16#153e# => read_data_o <= x"0000";
				when 16#153f# => read_data_o <= x"0000";
				when 16#1540# => read_data_o <= x"0000";
				when 16#1541# => read_data_o <= x"0000";
				when 16#1542# => read_data_o <= x"0000";
				when 16#1543# => read_data_o <= x"0000";
				when 16#1544# => read_data_o <= x"0000";
				when 16#1545# => read_data_o <= x"0000";
				when 16#1546# => read_data_o <= x"0000";
				when 16#1547# => read_data_o <= x"0000";
				when 16#1548# => read_data_o <= x"0000";
				when 16#1549# => read_data_o <= x"0000";
				when 16#154a# => read_data_o <= x"0000";
				when 16#154b# => read_data_o <= x"0000";
				when 16#154c# => read_data_o <= x"0000";
				when 16#154d# => read_data_o <= x"0000";
				when 16#154e# => read_data_o <= x"0000";
				when 16#154f# => read_data_o <= x"0000";
				when 16#1550# => read_data_o <= x"0000";
				when 16#1551# => read_data_o <= x"0000";
				when 16#1552# => read_data_o <= x"0000";
				when 16#1553# => read_data_o <= x"0000";
				when 16#1554# => read_data_o <= x"0000";
				when 16#1555# => read_data_o <= x"0000";
				when 16#1556# => read_data_o <= x"0000";
				when 16#1557# => read_data_o <= x"0000";
				when 16#1558# => read_data_o <= x"0000";
				when 16#1559# => read_data_o <= x"0000";
				when 16#155a# => read_data_o <= x"0000";
				when 16#155b# => read_data_o <= x"0000";
				when 16#155c# => read_data_o <= x"0000";
				when 16#155d# => read_data_o <= x"0000";
				when 16#155e# => read_data_o <= x"0000";
				when 16#155f# => read_data_o <= x"0000";
				when 16#1560# => read_data_o <= x"0000";
				when 16#1561# => read_data_o <= x"0000";
				when 16#1562# => read_data_o <= x"0000";
				when 16#1563# => read_data_o <= x"0000";
				when 16#1564# => read_data_o <= x"0000";
				when 16#1565# => read_data_o <= x"0000";
				when 16#1566# => read_data_o <= x"0000";
				when 16#1567# => read_data_o <= x"0000";
				when 16#1568# => read_data_o <= x"0000";
				when 16#1569# => read_data_o <= x"0000";
				when 16#156a# => read_data_o <= x"0000";
				when 16#156b# => read_data_o <= x"0000";
				when 16#156c# => read_data_o <= x"0000";
				when 16#156d# => read_data_o <= x"0000";
				when 16#156e# => read_data_o <= x"0000";
				when 16#156f# => read_data_o <= x"0000";
				when 16#1570# => read_data_o <= x"0000";
				when 16#1571# => read_data_o <= x"0000";
				when 16#1572# => read_data_o <= x"0000";
				when 16#1573# => read_data_o <= x"0000";
				when 16#1574# => read_data_o <= x"0000";
				when 16#1575# => read_data_o <= x"0000";
				when 16#1576# => read_data_o <= x"0000";
				when 16#1577# => read_data_o <= x"0000";
				when 16#1578# => read_data_o <= x"0000";
				when 16#1579# => read_data_o <= x"0000";
				when 16#157a# => read_data_o <= x"0000";
				when 16#157b# => read_data_o <= x"0000";
				when 16#157c# => read_data_o <= x"0000";
				when 16#157d# => read_data_o <= x"0000";
				when 16#157e# => read_data_o <= x"0000";
				when 16#157f# => read_data_o <= x"0000";
				when 16#1580# => read_data_o <= x"0000";
				when 16#1581# => read_data_o <= x"0000";
				when 16#1582# => read_data_o <= x"0000";
				when 16#1583# => read_data_o <= x"0000";
				when 16#1584# => read_data_o <= x"0000";
				when 16#1585# => read_data_o <= x"0000";
				when 16#1586# => read_data_o <= x"0000";
				when 16#1587# => read_data_o <= x"0000";
				when 16#1588# => read_data_o <= x"0000";
				when 16#1589# => read_data_o <= x"0000";
				when 16#158a# => read_data_o <= x"0000";
				when 16#158b# => read_data_o <= x"0000";
				when 16#158c# => read_data_o <= x"0000";
				when 16#158d# => read_data_o <= x"0000";
				when 16#158e# => read_data_o <= x"0000";
				when 16#158f# => read_data_o <= x"0000";
				when 16#1590# => read_data_o <= x"0000";
				when 16#1591# => read_data_o <= x"0000";
				when 16#1592# => read_data_o <= x"0000";
				when 16#1593# => read_data_o <= x"0000";
				when 16#1594# => read_data_o <= x"0000";
				when 16#1595# => read_data_o <= x"0000";
				when 16#1596# => read_data_o <= x"0000";
				when 16#1597# => read_data_o <= x"0000";
				when 16#1598# => read_data_o <= x"0000";
				when 16#1599# => read_data_o <= x"0000";
				when 16#159a# => read_data_o <= x"0000";
				when 16#159b# => read_data_o <= x"0000";
				when 16#159c# => read_data_o <= x"0000";
				when 16#159d# => read_data_o <= x"0000";
				when 16#159e# => read_data_o <= x"0000";
				when 16#159f# => read_data_o <= x"0000";
				when 16#15a0# => read_data_o <= x"0000";
				when 16#15a1# => read_data_o <= x"0000";
				when 16#15a2# => read_data_o <= x"0000";
				when 16#15a3# => read_data_o <= x"0000";
				when 16#15a4# => read_data_o <= x"0000";
				when 16#15a5# => read_data_o <= x"0000";
				when 16#15a6# => read_data_o <= x"0000";
				when 16#15a7# => read_data_o <= x"0000";
				when 16#15a8# => read_data_o <= x"0000";
				when 16#15a9# => read_data_o <= x"0000";
				when 16#15aa# => read_data_o <= x"0000";
				when 16#15ab# => read_data_o <= x"0000";
				when 16#15ac# => read_data_o <= x"0000";
				when 16#15ad# => read_data_o <= x"0000";
				when 16#15ae# => read_data_o <= x"0000";
				when 16#15af# => read_data_o <= x"0000";
				when 16#15b0# => read_data_o <= x"0000";
				when 16#15b1# => read_data_o <= x"0000";
				when 16#15b2# => read_data_o <= x"0000";
				when 16#15b3# => read_data_o <= x"0000";
				when 16#15b4# => read_data_o <= x"0000";
				when 16#15b5# => read_data_o <= x"0000";
				when 16#15b6# => read_data_o <= x"0000";
				when 16#15b7# => read_data_o <= x"0000";
				when 16#15b8# => read_data_o <= x"0000";
				when 16#15b9# => read_data_o <= x"0000";
				when 16#15ba# => read_data_o <= x"0000";
				when 16#15bb# => read_data_o <= x"0000";
				when 16#15bc# => read_data_o <= x"0000";
				when 16#15bd# => read_data_o <= x"0000";
				when 16#15be# => read_data_o <= x"0000";
				when 16#15bf# => read_data_o <= x"0000";
				when 16#15c0# => read_data_o <= x"0000";
				when 16#15c1# => read_data_o <= x"0000";
				when 16#15c2# => read_data_o <= x"0000";
				when 16#15c3# => read_data_o <= x"0000";
				when 16#15c4# => read_data_o <= x"0000";
				when 16#15c5# => read_data_o <= x"0000";
				when 16#15c6# => read_data_o <= x"0000";
				when 16#15c7# => read_data_o <= x"0000";
				when 16#15c8# => read_data_o <= x"0000";
				when 16#15c9# => read_data_o <= x"0000";
				when 16#15ca# => read_data_o <= x"0000";
				when 16#15cb# => read_data_o <= x"0000";
				when 16#15cc# => read_data_o <= x"0000";
				when 16#15cd# => read_data_o <= x"0000";
				when 16#15ce# => read_data_o <= x"0000";
				when 16#15cf# => read_data_o <= x"0000";
				when 16#15d0# => read_data_o <= x"0000";
				when 16#15d1# => read_data_o <= x"0000";
				when 16#15d2# => read_data_o <= x"0000";
				when 16#15d3# => read_data_o <= x"0000";
				when 16#15d4# => read_data_o <= x"0000";
				when 16#15d5# => read_data_o <= x"0000";
				when 16#15d6# => read_data_o <= x"0000";
				when 16#15d7# => read_data_o <= x"0000";
				when 16#15d8# => read_data_o <= x"0000";
				when 16#15d9# => read_data_o <= x"0000";
				when 16#15da# => read_data_o <= x"0000";
				when 16#15db# => read_data_o <= x"0000";
				when 16#15dc# => read_data_o <= x"0000";
				when 16#15dd# => read_data_o <= x"0000";
				when 16#15de# => read_data_o <= x"0000";
				when 16#15df# => read_data_o <= x"0000";
				when 16#15e0# => read_data_o <= x"0000";
				when 16#15e1# => read_data_o <= x"0000";
				when 16#15e2# => read_data_o <= x"0000";
				when 16#15e3# => read_data_o <= x"0000";
				when 16#15e4# => read_data_o <= x"0000";
				when 16#15e5# => read_data_o <= x"0000";
				when 16#15e6# => read_data_o <= x"0000";
				when 16#15e7# => read_data_o <= x"0000";
				when 16#15e8# => read_data_o <= x"0000";
				when 16#15e9# => read_data_o <= x"0000";
				when 16#15ea# => read_data_o <= x"0000";
				when 16#15eb# => read_data_o <= x"0000";
				when 16#15ec# => read_data_o <= x"0000";
				when 16#15ed# => read_data_o <= x"0000";
				when 16#15ee# => read_data_o <= x"0000";
				when 16#15ef# => read_data_o <= x"0000";
				when 16#15f0# => read_data_o <= x"0000";
				when 16#15f1# => read_data_o <= x"0000";
				when 16#15f2# => read_data_o <= x"0000";
				when 16#15f3# => read_data_o <= x"0000";
				when 16#15f4# => read_data_o <= x"0000";
				when 16#15f5# => read_data_o <= x"0000";
				when 16#15f6# => read_data_o <= x"0000";
				when 16#15f7# => read_data_o <= x"0000";
				when 16#15f8# => read_data_o <= x"0000";
				when 16#15f9# => read_data_o <= x"0000";
				when 16#15fa# => read_data_o <= x"0000";
				when 16#15fb# => read_data_o <= x"0000";
				when 16#15fc# => read_data_o <= x"0000";
				when 16#15fd# => read_data_o <= x"0000";
				when 16#15fe# => read_data_o <= x"0000";
				when 16#15ff# => read_data_o <= x"0000";
				when 16#1600# => read_data_o <= x"0000";
				when 16#1601# => read_data_o <= x"0000";
				when 16#1602# => read_data_o <= x"0000";
				when 16#1603# => read_data_o <= x"0000";
				when 16#1604# => read_data_o <= x"0000";
				when 16#1605# => read_data_o <= x"0000";
				when 16#1606# => read_data_o <= x"0000";
				when 16#1607# => read_data_o <= x"0000";
				when 16#1608# => read_data_o <= x"0000";
				when 16#1609# => read_data_o <= x"0000";
				when 16#160a# => read_data_o <= x"0000";
				when 16#160b# => read_data_o <= x"0000";
				when 16#160c# => read_data_o <= x"0000";
				when 16#160d# => read_data_o <= x"0000";
				when 16#160e# => read_data_o <= x"0000";
				when 16#160f# => read_data_o <= x"0000";
				when 16#1610# => read_data_o <= x"0000";
				when 16#1611# => read_data_o <= x"0000";
				when 16#1612# => read_data_o <= x"0000";
				when 16#1613# => read_data_o <= x"0000";
				when 16#1614# => read_data_o <= x"0000";
				when 16#1615# => read_data_o <= x"0000";
				when 16#1616# => read_data_o <= x"0000";
				when 16#1617# => read_data_o <= x"0000";
				when 16#1618# => read_data_o <= x"0000";
				when 16#1619# => read_data_o <= x"0000";
				when 16#161a# => read_data_o <= x"0000";
				when 16#161b# => read_data_o <= x"0000";
				when 16#161c# => read_data_o <= x"0000";
				when 16#161d# => read_data_o <= x"0000";
				when 16#161e# => read_data_o <= x"0000";
				when 16#161f# => read_data_o <= x"0000";
				when 16#1620# => read_data_o <= x"0000";
				when 16#1621# => read_data_o <= x"0000";
				when 16#1622# => read_data_o <= x"0000";
				when 16#1623# => read_data_o <= x"0000";
				when 16#1624# => read_data_o <= x"0000";
				when 16#1625# => read_data_o <= x"0000";
				when 16#1626# => read_data_o <= x"0000";
				when 16#1627# => read_data_o <= x"0000";
				when 16#1628# => read_data_o <= x"0000";
				when 16#1629# => read_data_o <= x"0000";
				when 16#162a# => read_data_o <= x"0000";
				when 16#162b# => read_data_o <= x"0000";
				when 16#162c# => read_data_o <= x"0000";
				when 16#162d# => read_data_o <= x"0000";
				when 16#162e# => read_data_o <= x"0000";
				when 16#162f# => read_data_o <= x"0000";
				when 16#1630# => read_data_o <= x"0000";
				when 16#1631# => read_data_o <= x"0000";
				when 16#1632# => read_data_o <= x"0000";
				when 16#1633# => read_data_o <= x"0000";
				when 16#1634# => read_data_o <= x"0000";
				when 16#1635# => read_data_o <= x"0000";
				when 16#1636# => read_data_o <= x"0000";
				when 16#1637# => read_data_o <= x"0000";
				when 16#1638# => read_data_o <= x"0000";
				when 16#1639# => read_data_o <= x"0000";
				when 16#163a# => read_data_o <= x"0000";
				when 16#163b# => read_data_o <= x"0000";
				when 16#163c# => read_data_o <= x"0000";
				when 16#163d# => read_data_o <= x"0000";
				when 16#163e# => read_data_o <= x"0000";
				when 16#163f# => read_data_o <= x"0000";
				when 16#1640# => read_data_o <= x"0000";
				when 16#1641# => read_data_o <= x"0000";
				when 16#1642# => read_data_o <= x"0000";
				when 16#1643# => read_data_o <= x"0000";
				when 16#1644# => read_data_o <= x"0000";
				when 16#1645# => read_data_o <= x"0000";
				when 16#1646# => read_data_o <= x"0000";
				when 16#1647# => read_data_o <= x"0000";
				when 16#1648# => read_data_o <= x"0000";
				when 16#1649# => read_data_o <= x"0000";
				when 16#164a# => read_data_o <= x"0000";
				when 16#164b# => read_data_o <= x"0000";
				when 16#164c# => read_data_o <= x"0000";
				when 16#164d# => read_data_o <= x"0000";
				when 16#164e# => read_data_o <= x"0000";
				when 16#164f# => read_data_o <= x"0000";
				when 16#1650# => read_data_o <= x"0000";
				when 16#1651# => read_data_o <= x"0000";
				when 16#1652# => read_data_o <= x"0000";
				when 16#1653# => read_data_o <= x"0000";
				when 16#1654# => read_data_o <= x"0000";
				when 16#1655# => read_data_o <= x"0000";
				when 16#1656# => read_data_o <= x"0000";
				when 16#1657# => read_data_o <= x"0000";
				when 16#1658# => read_data_o <= x"0000";
				when 16#1659# => read_data_o <= x"0000";
				when 16#165a# => read_data_o <= x"0000";
				when 16#165b# => read_data_o <= x"0000";
				when 16#165c# => read_data_o <= x"0000";
				when 16#165d# => read_data_o <= x"0000";
				when 16#165e# => read_data_o <= x"0000";
				when 16#165f# => read_data_o <= x"0000";
				when 16#1660# => read_data_o <= x"0000";
				when 16#1661# => read_data_o <= x"0000";
				when 16#1662# => read_data_o <= x"0000";
				when 16#1663# => read_data_o <= x"0000";
				when 16#1664# => read_data_o <= x"0000";
				when 16#1665# => read_data_o <= x"0000";
				when 16#1666# => read_data_o <= x"0000";
				when 16#1667# => read_data_o <= x"0000";
				when 16#1668# => read_data_o <= x"0000";
				when 16#1669# => read_data_o <= x"0000";
				when 16#166a# => read_data_o <= x"0000";
				when 16#166b# => read_data_o <= x"0000";
				when 16#166c# => read_data_o <= x"0000";
				when 16#166d# => read_data_o <= x"0000";
				when 16#166e# => read_data_o <= x"0000";
				when 16#166f# => read_data_o <= x"0000";
				when 16#1670# => read_data_o <= x"0000";
				when 16#1671# => read_data_o <= x"0000";
				when 16#1672# => read_data_o <= x"0000";
				when 16#1673# => read_data_o <= x"0000";
				when 16#1674# => read_data_o <= x"0000";
				when 16#1675# => read_data_o <= x"0000";
				when 16#1676# => read_data_o <= x"0000";
				when 16#1677# => read_data_o <= x"0000";
				when 16#1678# => read_data_o <= x"0000";
				when 16#1679# => read_data_o <= x"0000";
				when 16#167a# => read_data_o <= x"0000";
				when 16#167b# => read_data_o <= x"0000";
				when 16#167c# => read_data_o <= x"0000";
				when 16#167d# => read_data_o <= x"0000";
				when 16#167e# => read_data_o <= x"0000";
				when 16#167f# => read_data_o <= x"0000";
				when 16#1680# => read_data_o <= x"0000";
				when 16#1681# => read_data_o <= x"0000";
				when 16#1682# => read_data_o <= x"0000";
				when 16#1683# => read_data_o <= x"0000";
				when 16#1684# => read_data_o <= x"0000";
				when 16#1685# => read_data_o <= x"0000";
				when 16#1686# => read_data_o <= x"0000";
				when 16#1687# => read_data_o <= x"0000";
				when 16#1688# => read_data_o <= x"0000";
				when 16#1689# => read_data_o <= x"0000";
				when 16#168a# => read_data_o <= x"0000";
				when 16#168b# => read_data_o <= x"0000";
				when 16#168c# => read_data_o <= x"0000";
				when 16#168d# => read_data_o <= x"0000";
				when 16#168e# => read_data_o <= x"0000";
				when 16#168f# => read_data_o <= x"0000";
				when 16#1690# => read_data_o <= x"0000";
				when 16#1691# => read_data_o <= x"0000";
				when 16#1692# => read_data_o <= x"0000";
				when 16#1693# => read_data_o <= x"0000";
				when 16#1694# => read_data_o <= x"0000";
				when 16#1695# => read_data_o <= x"0000";
				when 16#1696# => read_data_o <= x"0000";
				when 16#1697# => read_data_o <= x"0000";
				when 16#1698# => read_data_o <= x"0000";
				when 16#1699# => read_data_o <= x"0000";
				when 16#169a# => read_data_o <= x"0000";
				when 16#169b# => read_data_o <= x"0000";
				when 16#169c# => read_data_o <= x"0000";
				when 16#169d# => read_data_o <= x"0000";
				when 16#169e# => read_data_o <= x"0000";
				when 16#169f# => read_data_o <= x"0000";
				when 16#16a0# => read_data_o <= x"0000";
				when 16#16a1# => read_data_o <= x"0000";
				when 16#16a2# => read_data_o <= x"0000";
				when 16#16a3# => read_data_o <= x"0000";
				when 16#16a4# => read_data_o <= x"0000";
				when 16#16a5# => read_data_o <= x"0000";
				when 16#16a6# => read_data_o <= x"0000";
				when 16#16a7# => read_data_o <= x"0000";
				when 16#16a8# => read_data_o <= x"0000";
				when 16#16a9# => read_data_o <= x"0000";
				when 16#16aa# => read_data_o <= x"0000";
				when 16#16ab# => read_data_o <= x"0000";
				when 16#16ac# => read_data_o <= x"0000";
				when 16#16ad# => read_data_o <= x"0000";
				when 16#16ae# => read_data_o <= x"0000";
				when 16#16af# => read_data_o <= x"0000";
				when 16#16b0# => read_data_o <= x"0000";
				when 16#16b1# => read_data_o <= x"0000";
				when 16#16b2# => read_data_o <= x"0000";
				when 16#16b3# => read_data_o <= x"0000";
				when 16#16b4# => read_data_o <= x"0000";
				when 16#16b5# => read_data_o <= x"0000";
				when 16#16b6# => read_data_o <= x"0000";
				when 16#16b7# => read_data_o <= x"0000";
				when 16#16b8# => read_data_o <= x"0000";
				when 16#16b9# => read_data_o <= x"0000";
				when 16#16ba# => read_data_o <= x"0000";
				when 16#16bb# => read_data_o <= x"0000";
				when 16#16bc# => read_data_o <= x"0000";
				when 16#16bd# => read_data_o <= x"0000";
				when 16#16be# => read_data_o <= x"0000";
				when 16#16bf# => read_data_o <= x"0000";
				when 16#16c0# => read_data_o <= x"0000";
				when 16#16c1# => read_data_o <= x"0000";
				when 16#16c2# => read_data_o <= x"0000";
				when 16#16c3# => read_data_o <= x"0000";
				when 16#16c4# => read_data_o <= x"0000";
				when 16#16c5# => read_data_o <= x"0000";
				when 16#16c6# => read_data_o <= x"0000";
				when 16#16c7# => read_data_o <= x"0000";
				when 16#16c8# => read_data_o <= x"0000";
				when 16#16c9# => read_data_o <= x"0000";
				when 16#16ca# => read_data_o <= x"0000";
				when 16#16cb# => read_data_o <= x"0000";
				when 16#16cc# => read_data_o <= x"0000";
				when 16#16cd# => read_data_o <= x"0000";
				when 16#16ce# => read_data_o <= x"0000";
				when 16#16cf# => read_data_o <= x"0000";
				when 16#16d0# => read_data_o <= x"0000";
				when 16#16d1# => read_data_o <= x"0000";
				when 16#16d2# => read_data_o <= x"0000";
				when 16#16d3# => read_data_o <= x"0000";
				when 16#16d4# => read_data_o <= x"0000";
				when 16#16d5# => read_data_o <= x"0000";
				when 16#16d6# => read_data_o <= x"0000";
				when 16#16d7# => read_data_o <= x"0000";
				when 16#16d8# => read_data_o <= x"0000";
				when 16#16d9# => read_data_o <= x"0000";
				when 16#16da# => read_data_o <= x"0000";
				when 16#16db# => read_data_o <= x"0000";
				when 16#16dc# => read_data_o <= x"0000";
				when 16#16dd# => read_data_o <= x"0000";
				when 16#16de# => read_data_o <= x"0000";
				when 16#16df# => read_data_o <= x"0000";
				when 16#16e0# => read_data_o <= x"0000";
				when 16#16e1# => read_data_o <= x"0000";
				when 16#16e2# => read_data_o <= x"0000";
				when 16#16e3# => read_data_o <= x"0000";
				when 16#16e4# => read_data_o <= x"0000";
				when 16#16e5# => read_data_o <= x"0000";
				when 16#16e6# => read_data_o <= x"0000";
				when 16#16e7# => read_data_o <= x"0000";
				when 16#16e8# => read_data_o <= x"0000";
				when 16#16e9# => read_data_o <= x"0000";
				when 16#16ea# => read_data_o <= x"0000";
				when 16#16eb# => read_data_o <= x"0000";
				when 16#16ec# => read_data_o <= x"0000";
				when 16#16ed# => read_data_o <= x"0000";
				when 16#16ee# => read_data_o <= x"0000";
				when 16#16ef# => read_data_o <= x"0000";
				when 16#16f0# => read_data_o <= x"0000";
				when 16#16f1# => read_data_o <= x"0000";
				when 16#16f2# => read_data_o <= x"0000";
				when 16#16f3# => read_data_o <= x"0000";
				when 16#16f4# => read_data_o <= x"0000";
				when 16#16f5# => read_data_o <= x"0000";
				when 16#16f6# => read_data_o <= x"0000";
				when 16#16f7# => read_data_o <= x"0000";
				when 16#16f8# => read_data_o <= x"0000";
				when 16#16f9# => read_data_o <= x"0000";
				when 16#16fa# => read_data_o <= x"0000";
				when 16#16fb# => read_data_o <= x"0000";
				when 16#16fc# => read_data_o <= x"0000";
				when 16#16fd# => read_data_o <= x"0000";
				when 16#16fe# => read_data_o <= x"0000";
				when 16#16ff# => read_data_o <= x"0000";
				when 16#1700# => read_data_o <= x"0000";
				when 16#1701# => read_data_o <= x"0000";
				when 16#1702# => read_data_o <= x"0000";
				when 16#1703# => read_data_o <= x"0000";
				when 16#1704# => read_data_o <= x"0000";
				when 16#1705# => read_data_o <= x"0000";
				when 16#1706# => read_data_o <= x"0000";
				when 16#1707# => read_data_o <= x"0000";
				when 16#1708# => read_data_o <= x"0000";
				when 16#1709# => read_data_o <= x"0000";
				when 16#170a# => read_data_o <= x"0000";
				when 16#170b# => read_data_o <= x"0000";
				when 16#170c# => read_data_o <= x"0000";
				when 16#170d# => read_data_o <= x"0000";
				when 16#170e# => read_data_o <= x"0000";
				when 16#170f# => read_data_o <= x"0000";
				when 16#1710# => read_data_o <= x"0000";
				when 16#1711# => read_data_o <= x"0000";
				when 16#1712# => read_data_o <= x"0000";
				when 16#1713# => read_data_o <= x"0000";
				when 16#1714# => read_data_o <= x"0000";
				when 16#1715# => read_data_o <= x"0000";
				when 16#1716# => read_data_o <= x"0000";
				when 16#1717# => read_data_o <= x"0000";
				when 16#1718# => read_data_o <= x"0000";
				when 16#1719# => read_data_o <= x"0000";
				when 16#171a# => read_data_o <= x"0000";
				when 16#171b# => read_data_o <= x"0000";
				when 16#171c# => read_data_o <= x"0000";
				when 16#171d# => read_data_o <= x"0000";
				when 16#171e# => read_data_o <= x"0000";
				when 16#171f# => read_data_o <= x"0000";
				when 16#1720# => read_data_o <= x"0000";
				when 16#1721# => read_data_o <= x"0000";
				when 16#1722# => read_data_o <= x"0000";
				when 16#1723# => read_data_o <= x"0000";
				when 16#1724# => read_data_o <= x"0000";
				when 16#1725# => read_data_o <= x"0000";
				when 16#1726# => read_data_o <= x"0000";
				when 16#1727# => read_data_o <= x"0000";
				when 16#1728# => read_data_o <= x"0000";
				when 16#1729# => read_data_o <= x"0000";
				when 16#172a# => read_data_o <= x"0000";
				when 16#172b# => read_data_o <= x"0000";
				when 16#172c# => read_data_o <= x"0000";
				when 16#172d# => read_data_o <= x"0000";
				when 16#172e# => read_data_o <= x"0000";
				when 16#172f# => read_data_o <= x"0000";
				when 16#1730# => read_data_o <= x"0000";
				when 16#1731# => read_data_o <= x"0000";
				when 16#1732# => read_data_o <= x"0000";
				when 16#1733# => read_data_o <= x"0000";
				when 16#1734# => read_data_o <= x"0000";
				when 16#1735# => read_data_o <= x"0000";
				when 16#1736# => read_data_o <= x"0000";
				when 16#1737# => read_data_o <= x"0000";
				when 16#1738# => read_data_o <= x"0000";
				when 16#1739# => read_data_o <= x"0000";
				when 16#173a# => read_data_o <= x"0000";
				when 16#173b# => read_data_o <= x"0000";
				when 16#173c# => read_data_o <= x"0000";
				when 16#173d# => read_data_o <= x"0000";
				when 16#173e# => read_data_o <= x"0000";
				when 16#173f# => read_data_o <= x"0000";
				when 16#1740# => read_data_o <= x"0000";
				when 16#1741# => read_data_o <= x"0000";
				when 16#1742# => read_data_o <= x"0000";
				when 16#1743# => read_data_o <= x"0000";
				when 16#1744# => read_data_o <= x"0000";
				when 16#1745# => read_data_o <= x"0000";
				when 16#1746# => read_data_o <= x"0000";
				when 16#1747# => read_data_o <= x"0000";
				when 16#1748# => read_data_o <= x"0000";
				when 16#1749# => read_data_o <= x"0000";
				when 16#174a# => read_data_o <= x"0000";
				when 16#174b# => read_data_o <= x"0000";
				when 16#174c# => read_data_o <= x"0000";
				when 16#174d# => read_data_o <= x"0000";
				when 16#174e# => read_data_o <= x"0000";
				when 16#174f# => read_data_o <= x"0000";
				when 16#1750# => read_data_o <= x"0000";
				when 16#1751# => read_data_o <= x"0000";
				when 16#1752# => read_data_o <= x"0000";
				when 16#1753# => read_data_o <= x"0000";
				when 16#1754# => read_data_o <= x"0000";
				when 16#1755# => read_data_o <= x"0000";
				when 16#1756# => read_data_o <= x"0000";
				when 16#1757# => read_data_o <= x"0000";
				when 16#1758# => read_data_o <= x"0000";
				when 16#1759# => read_data_o <= x"0000";
				when 16#175a# => read_data_o <= x"0000";
				when 16#175b# => read_data_o <= x"0000";
				when 16#175c# => read_data_o <= x"0000";
				when 16#175d# => read_data_o <= x"0000";
				when 16#175e# => read_data_o <= x"0000";
				when 16#175f# => read_data_o <= x"0000";
				when 16#1760# => read_data_o <= x"0000";
				when 16#1761# => read_data_o <= x"0000";
				when 16#1762# => read_data_o <= x"0000";
				when 16#1763# => read_data_o <= x"0000";
				when 16#1764# => read_data_o <= x"0000";
				when 16#1765# => read_data_o <= x"0000";
				when 16#1766# => read_data_o <= x"0000";
				when 16#1767# => read_data_o <= x"0000";
				when 16#1768# => read_data_o <= x"0000";
				when 16#1769# => read_data_o <= x"0000";
				when 16#176a# => read_data_o <= x"0000";
				when 16#176b# => read_data_o <= x"0000";
				when 16#176c# => read_data_o <= x"0000";
				when 16#176d# => read_data_o <= x"0000";
				when 16#176e# => read_data_o <= x"0000";
				when 16#176f# => read_data_o <= x"0000";
				when 16#1770# => read_data_o <= x"0000";
				when 16#1771# => read_data_o <= x"0000";
				when 16#1772# => read_data_o <= x"0000";
				when 16#1773# => read_data_o <= x"0000";
				when 16#1774# => read_data_o <= x"0000";
				when 16#1775# => read_data_o <= x"0000";
				when 16#1776# => read_data_o <= x"0000";
				when 16#1777# => read_data_o <= x"0000";
				when 16#1778# => read_data_o <= x"0000";
				when 16#1779# => read_data_o <= x"0000";
				when 16#177a# => read_data_o <= x"0000";
				when 16#177b# => read_data_o <= x"0000";
				when 16#177c# => read_data_o <= x"0000";
				when 16#177d# => read_data_o <= x"0000";
				when 16#177e# => read_data_o <= x"0000";
				when 16#177f# => read_data_o <= x"0000";
				when 16#1780# => read_data_o <= x"0000";
				when 16#1781# => read_data_o <= x"0000";
				when 16#1782# => read_data_o <= x"0000";
				when 16#1783# => read_data_o <= x"0000";
				when 16#1784# => read_data_o <= x"0000";
				when 16#1785# => read_data_o <= x"0000";
				when 16#1786# => read_data_o <= x"0000";
				when 16#1787# => read_data_o <= x"0000";
				when 16#1788# => read_data_o <= x"0000";
				when 16#1789# => read_data_o <= x"0000";
				when 16#178a# => read_data_o <= x"0000";
				when 16#178b# => read_data_o <= x"0000";
				when 16#178c# => read_data_o <= x"0000";
				when 16#178d# => read_data_o <= x"0000";
				when 16#178e# => read_data_o <= x"0000";
				when 16#178f# => read_data_o <= x"0000";
				when 16#1790# => read_data_o <= x"0000";
				when 16#1791# => read_data_o <= x"0000";
				when 16#1792# => read_data_o <= x"0000";
				when 16#1793# => read_data_o <= x"0000";
				when 16#1794# => read_data_o <= x"0000";
				when 16#1795# => read_data_o <= x"0000";
				when 16#1796# => read_data_o <= x"0000";
				when 16#1797# => read_data_o <= x"0000";
				when 16#1798# => read_data_o <= x"0000";
				when 16#1799# => read_data_o <= x"0000";
				when 16#179a# => read_data_o <= x"0000";
				when 16#179b# => read_data_o <= x"0000";
				when 16#179c# => read_data_o <= x"0000";
				when 16#179d# => read_data_o <= x"0000";
				when 16#179e# => read_data_o <= x"0000";
				when 16#179f# => read_data_o <= x"0000";
				when 16#17a0# => read_data_o <= x"0000";
				when 16#17a1# => read_data_o <= x"0000";
				when 16#17a2# => read_data_o <= x"0000";
				when 16#17a3# => read_data_o <= x"0000";
				when 16#17a4# => read_data_o <= x"0000";
				when 16#17a5# => read_data_o <= x"0000";
				when 16#17a6# => read_data_o <= x"0000";
				when 16#17a7# => read_data_o <= x"0000";
				when 16#17a8# => read_data_o <= x"0000";
				when 16#17a9# => read_data_o <= x"0000";
				when 16#17aa# => read_data_o <= x"0000";
				when 16#17ab# => read_data_o <= x"0000";
				when 16#17ac# => read_data_o <= x"0000";
				when 16#17ad# => read_data_o <= x"0000";
				when 16#17ae# => read_data_o <= x"0000";
				when 16#17af# => read_data_o <= x"0000";
				when 16#17b0# => read_data_o <= x"0000";
				when 16#17b1# => read_data_o <= x"0000";
				when 16#17b2# => read_data_o <= x"0000";
				when 16#17b3# => read_data_o <= x"0000";
				when 16#17b4# => read_data_o <= x"0000";
				when 16#17b5# => read_data_o <= x"0000";
				when 16#17b6# => read_data_o <= x"0000";
				when 16#17b7# => read_data_o <= x"0000";
				when 16#17b8# => read_data_o <= x"0000";
				when 16#17b9# => read_data_o <= x"0000";
				when 16#17ba# => read_data_o <= x"0000";
				when 16#17bb# => read_data_o <= x"0000";
				when 16#17bc# => read_data_o <= x"0000";
				when 16#17bd# => read_data_o <= x"0000";
				when 16#17be# => read_data_o <= x"0000";
				when 16#17bf# => read_data_o <= x"0000";
				when 16#17c0# => read_data_o <= x"0000";
				when 16#17c1# => read_data_o <= x"0000";
				when 16#17c2# => read_data_o <= x"0000";
				when 16#17c3# => read_data_o <= x"0000";
				when 16#17c4# => read_data_o <= x"0000";
				when 16#17c5# => read_data_o <= x"0000";
				when 16#17c6# => read_data_o <= x"0000";
				when 16#17c7# => read_data_o <= x"0000";
				when 16#17c8# => read_data_o <= x"0000";
				when 16#17c9# => read_data_o <= x"0000";
				when 16#17ca# => read_data_o <= x"0000";
				when 16#17cb# => read_data_o <= x"0000";
				when 16#17cc# => read_data_o <= x"0000";
				when 16#17cd# => read_data_o <= x"0000";
				when 16#17ce# => read_data_o <= x"0000";
				when 16#17cf# => read_data_o <= x"0000";
				when 16#17d0# => read_data_o <= x"0000";
				when 16#17d1# => read_data_o <= x"0000";
				when 16#17d2# => read_data_o <= x"0000";
				when 16#17d3# => read_data_o <= x"0000";
				when 16#17d4# => read_data_o <= x"0000";
				when 16#17d5# => read_data_o <= x"0000";
				when 16#17d6# => read_data_o <= x"0000";
				when 16#17d7# => read_data_o <= x"0000";
				when 16#17d8# => read_data_o <= x"0000";
				when 16#17d9# => read_data_o <= x"0000";
				when 16#17da# => read_data_o <= x"0000";
				when 16#17db# => read_data_o <= x"0000";
				when 16#17dc# => read_data_o <= x"0000";
				when 16#17dd# => read_data_o <= x"0000";
				when 16#17de# => read_data_o <= x"0000";
				when 16#17df# => read_data_o <= x"0000";
				when 16#17e0# => read_data_o <= x"0000";
				when 16#17e1# => read_data_o <= x"0000";
				when 16#17e2# => read_data_o <= x"0000";
				when 16#17e3# => read_data_o <= x"0000";
				when 16#17e4# => read_data_o <= x"0000";
				when 16#17e5# => read_data_o <= x"0000";
				when 16#17e6# => read_data_o <= x"0000";
				when 16#17e7# => read_data_o <= x"0000";
				when 16#17e8# => read_data_o <= x"0000";
				when 16#17e9# => read_data_o <= x"0000";
				when 16#17ea# => read_data_o <= x"0000";
				when 16#17eb# => read_data_o <= x"0000";
				when 16#17ec# => read_data_o <= x"0000";
				when 16#17ed# => read_data_o <= x"0000";
				when 16#17ee# => read_data_o <= x"0000";
				when 16#17ef# => read_data_o <= x"0000";
				when 16#17f0# => read_data_o <= x"0000";
				when 16#17f1# => read_data_o <= x"0000";
				when 16#17f2# => read_data_o <= x"0000";
				when 16#17f3# => read_data_o <= x"0000";
				when 16#17f4# => read_data_o <= x"0000";
				when 16#17f5# => read_data_o <= x"0000";
				when 16#17f6# => read_data_o <= x"0000";
				when 16#17f7# => read_data_o <= x"0000";
				when 16#17f8# => read_data_o <= x"0000";
				when 16#17f9# => read_data_o <= x"0000";
				when 16#17fa# => read_data_o <= x"0000";
				when 16#17fb# => read_data_o <= x"0000";
				when 16#17fc# => read_data_o <= x"0000";
				when 16#17fd# => read_data_o <= x"0000";
				when 16#17fe# => read_data_o <= x"0000";
				when 16#17ff# => read_data_o <= x"0000";
				when 16#1800# => read_data_o <= x"0000";
				when 16#1801# => read_data_o <= x"0000";
				when 16#1802# => read_data_o <= x"0000";
				when 16#1803# => read_data_o <= x"0000";
				when 16#1804# => read_data_o <= x"0000";
				when 16#1805# => read_data_o <= x"0000";
				when 16#1806# => read_data_o <= x"0000";
				when 16#1807# => read_data_o <= x"0000";
				when 16#1808# => read_data_o <= x"0000";
				when 16#1809# => read_data_o <= x"0000";
				when 16#180a# => read_data_o <= x"0000";
				when 16#180b# => read_data_o <= x"0000";
				when 16#180c# => read_data_o <= x"0000";
				when 16#180d# => read_data_o <= x"0000";
				when 16#180e# => read_data_o <= x"0000";
				when 16#180f# => read_data_o <= x"0000";
				when 16#1810# => read_data_o <= x"0000";
				when 16#1811# => read_data_o <= x"0000";
				when 16#1812# => read_data_o <= x"0000";
				when 16#1813# => read_data_o <= x"0000";
				when 16#1814# => read_data_o <= x"0000";
				when 16#1815# => read_data_o <= x"0000";
				when 16#1816# => read_data_o <= x"0000";
				when 16#1817# => read_data_o <= x"0000";
				when 16#1818# => read_data_o <= x"0000";
				when 16#1819# => read_data_o <= x"0000";
				when 16#181a# => read_data_o <= x"0000";
				when 16#181b# => read_data_o <= x"0000";
				when 16#181c# => read_data_o <= x"0000";
				when 16#181d# => read_data_o <= x"0000";
				when 16#181e# => read_data_o <= x"0000";
				when 16#181f# => read_data_o <= x"0000";
				when 16#1820# => read_data_o <= x"0000";
				when 16#1821# => read_data_o <= x"0000";
				when 16#1822# => read_data_o <= x"0000";
				when 16#1823# => read_data_o <= x"0000";
				when 16#1824# => read_data_o <= x"0000";
				when 16#1825# => read_data_o <= x"0000";
				when 16#1826# => read_data_o <= x"0000";
				when 16#1827# => read_data_o <= x"0000";
				when 16#1828# => read_data_o <= x"0000";
				when 16#1829# => read_data_o <= x"0000";
				when 16#182a# => read_data_o <= x"0000";
				when 16#182b# => read_data_o <= x"0000";
				when 16#182c# => read_data_o <= x"0000";
				when 16#182d# => read_data_o <= x"0000";
				when 16#182e# => read_data_o <= x"0000";
				when 16#182f# => read_data_o <= x"0000";
				when 16#1830# => read_data_o <= x"0000";
				when 16#1831# => read_data_o <= x"0000";
				when 16#1832# => read_data_o <= x"0000";
				when 16#1833# => read_data_o <= x"0000";
				when 16#1834# => read_data_o <= x"0000";
				when 16#1835# => read_data_o <= x"0000";
				when 16#1836# => read_data_o <= x"0000";
				when 16#1837# => read_data_o <= x"0000";
				when 16#1838# => read_data_o <= x"0000";
				when 16#1839# => read_data_o <= x"0000";
				when 16#183a# => read_data_o <= x"0000";
				when 16#183b# => read_data_o <= x"0000";
				when 16#183c# => read_data_o <= x"0000";
				when 16#183d# => read_data_o <= x"0000";
				when 16#183e# => read_data_o <= x"0000";
				when 16#183f# => read_data_o <= x"0000";
				when 16#1840# => read_data_o <= x"0000";
				when 16#1841# => read_data_o <= x"0000";
				when 16#1842# => read_data_o <= x"0000";
				when 16#1843# => read_data_o <= x"0000";
				when 16#1844# => read_data_o <= x"0000";
				when 16#1845# => read_data_o <= x"0000";
				when 16#1846# => read_data_o <= x"0000";
				when 16#1847# => read_data_o <= x"0000";
				when 16#1848# => read_data_o <= x"0000";
				when 16#1849# => read_data_o <= x"0000";
				when 16#184a# => read_data_o <= x"0000";
				when 16#184b# => read_data_o <= x"0000";
				when 16#184c# => read_data_o <= x"0000";
				when 16#184d# => read_data_o <= x"0000";
				when 16#184e# => read_data_o <= x"0000";
				when 16#184f# => read_data_o <= x"0000";
				when 16#1850# => read_data_o <= x"0000";
				when 16#1851# => read_data_o <= x"0000";
				when 16#1852# => read_data_o <= x"0000";
				when 16#1853# => read_data_o <= x"0000";
				when 16#1854# => read_data_o <= x"0000";
				when 16#1855# => read_data_o <= x"0000";
				when 16#1856# => read_data_o <= x"0000";
				when 16#1857# => read_data_o <= x"0000";
				when 16#1858# => read_data_o <= x"0000";
				when 16#1859# => read_data_o <= x"0000";
				when 16#185a# => read_data_o <= x"0000";
				when 16#185b# => read_data_o <= x"0000";
				when 16#185c# => read_data_o <= x"0000";
				when 16#185d# => read_data_o <= x"0000";
				when 16#185e# => read_data_o <= x"0000";
				when 16#185f# => read_data_o <= x"0000";
				when 16#1860# => read_data_o <= x"0000";
				when 16#1861# => read_data_o <= x"0000";
				when 16#1862# => read_data_o <= x"0000";
				when 16#1863# => read_data_o <= x"0000";
				when 16#1864# => read_data_o <= x"0000";
				when 16#1865# => read_data_o <= x"0000";
				when 16#1866# => read_data_o <= x"0000";
				when 16#1867# => read_data_o <= x"0000";
				when 16#1868# => read_data_o <= x"0000";
				when 16#1869# => read_data_o <= x"0000";
				when 16#186a# => read_data_o <= x"0000";
				when 16#186b# => read_data_o <= x"0000";
				when 16#186c# => read_data_o <= x"0000";
				when 16#186d# => read_data_o <= x"0000";
				when 16#186e# => read_data_o <= x"0000";
				when 16#186f# => read_data_o <= x"0000";
				when 16#1870# => read_data_o <= x"0000";
				when 16#1871# => read_data_o <= x"0000";
				when 16#1872# => read_data_o <= x"0000";
				when 16#1873# => read_data_o <= x"0000";
				when 16#1874# => read_data_o <= x"0000";
				when 16#1875# => read_data_o <= x"0000";
				when 16#1876# => read_data_o <= x"0000";
				when 16#1877# => read_data_o <= x"0000";
				when 16#1878# => read_data_o <= x"0000";
				when 16#1879# => read_data_o <= x"0000";
				when 16#187a# => read_data_o <= x"0000";
				when 16#187b# => read_data_o <= x"0000";
				when 16#187c# => read_data_o <= x"0000";
				when 16#187d# => read_data_o <= x"0000";
				when 16#187e# => read_data_o <= x"0000";
				when 16#187f# => read_data_o <= x"0000";
				when 16#1880# => read_data_o <= x"0000";
				when 16#1881# => read_data_o <= x"0000";
				when 16#1882# => read_data_o <= x"0000";
				when 16#1883# => read_data_o <= x"0000";
				when 16#1884# => read_data_o <= x"0000";
				when 16#1885# => read_data_o <= x"0000";
				when 16#1886# => read_data_o <= x"0000";
				when 16#1887# => read_data_o <= x"0000";
				when 16#1888# => read_data_o <= x"0000";
				when 16#1889# => read_data_o <= x"0000";
				when 16#188a# => read_data_o <= x"0000";
				when 16#188b# => read_data_o <= x"0000";
				when 16#188c# => read_data_o <= x"0000";
				when 16#188d# => read_data_o <= x"0000";
				when 16#188e# => read_data_o <= x"0000";
				when 16#188f# => read_data_o <= x"0000";
				when 16#1890# => read_data_o <= x"0000";
				when 16#1891# => read_data_o <= x"0000";
				when 16#1892# => read_data_o <= x"0000";
				when 16#1893# => read_data_o <= x"0000";
				when 16#1894# => read_data_o <= x"0000";
				when 16#1895# => read_data_o <= x"0000";
				when 16#1896# => read_data_o <= x"0000";
				when 16#1897# => read_data_o <= x"0000";
				when 16#1898# => read_data_o <= x"0000";
				when 16#1899# => read_data_o <= x"0000";
				when 16#189a# => read_data_o <= x"0000";
				when 16#189b# => read_data_o <= x"0000";
				when 16#189c# => read_data_o <= x"0000";
				when 16#189d# => read_data_o <= x"0000";
				when 16#189e# => read_data_o <= x"0000";
				when 16#189f# => read_data_o <= x"0000";
				when 16#18a0# => read_data_o <= x"0000";
				when 16#18a1# => read_data_o <= x"0000";
				when 16#18a2# => read_data_o <= x"0000";
				when 16#18a3# => read_data_o <= x"0000";
				when 16#18a4# => read_data_o <= x"0000";
				when 16#18a5# => read_data_o <= x"0000";
				when 16#18a6# => read_data_o <= x"0000";
				when 16#18a7# => read_data_o <= x"0000";
				when 16#18a8# => read_data_o <= x"0000";
				when 16#18a9# => read_data_o <= x"0000";
				when 16#18aa# => read_data_o <= x"0000";
				when 16#18ab# => read_data_o <= x"0000";
				when 16#18ac# => read_data_o <= x"0000";
				when 16#18ad# => read_data_o <= x"0000";
				when 16#18ae# => read_data_o <= x"0000";
				when 16#18af# => read_data_o <= x"0000";
				when 16#18b0# => read_data_o <= x"0000";
				when 16#18b1# => read_data_o <= x"0000";
				when 16#18b2# => read_data_o <= x"0000";
				when 16#18b3# => read_data_o <= x"0000";
				when 16#18b4# => read_data_o <= x"0000";
				when 16#18b5# => read_data_o <= x"0000";
				when 16#18b6# => read_data_o <= x"0000";
				when 16#18b7# => read_data_o <= x"0000";
				when 16#18b8# => read_data_o <= x"0000";
				when 16#18b9# => read_data_o <= x"0000";
				when 16#18ba# => read_data_o <= x"0000";
				when 16#18bb# => read_data_o <= x"0000";
				when 16#18bc# => read_data_o <= x"0000";
				when 16#18bd# => read_data_o <= x"0000";
				when 16#18be# => read_data_o <= x"0000";
				when 16#18bf# => read_data_o <= x"0000";
				when 16#18c0# => read_data_o <= x"0000";
				when 16#18c1# => read_data_o <= x"0000";
				when 16#18c2# => read_data_o <= x"0000";
				when 16#18c3# => read_data_o <= x"0000";
				when 16#18c4# => read_data_o <= x"0000";
				when 16#18c5# => read_data_o <= x"0000";
				when 16#18c6# => read_data_o <= x"0000";
				when 16#18c7# => read_data_o <= x"0000";
				when 16#18c8# => read_data_o <= x"0000";
				when 16#18c9# => read_data_o <= x"0000";
				when 16#18ca# => read_data_o <= x"0000";
				when 16#18cb# => read_data_o <= x"0000";
				when 16#18cc# => read_data_o <= x"0000";
				when 16#18cd# => read_data_o <= x"0000";
				when 16#18ce# => read_data_o <= x"0000";
				when 16#18cf# => read_data_o <= x"0000";
				when 16#18d0# => read_data_o <= x"0000";
				when 16#18d1# => read_data_o <= x"0000";
				when 16#18d2# => read_data_o <= x"0000";
				when 16#18d3# => read_data_o <= x"0000";
				when 16#18d4# => read_data_o <= x"0000";
				when 16#18d5# => read_data_o <= x"0000";
				when 16#18d6# => read_data_o <= x"0000";
				when 16#18d7# => read_data_o <= x"0000";
				when 16#18d8# => read_data_o <= x"0000";
				when 16#18d9# => read_data_o <= x"0000";
				when 16#18da# => read_data_o <= x"0000";
				when 16#18db# => read_data_o <= x"0000";
				when 16#18dc# => read_data_o <= x"0000";
				when 16#18dd# => read_data_o <= x"0000";
				when 16#18de# => read_data_o <= x"0000";
				when 16#18df# => read_data_o <= x"0000";
				when 16#18e0# => read_data_o <= x"0000";
				when 16#18e1# => read_data_o <= x"0000";
				when 16#18e2# => read_data_o <= x"0000";
				when 16#18e3# => read_data_o <= x"0000";
				when 16#18e4# => read_data_o <= x"0000";
				when 16#18e5# => read_data_o <= x"0000";
				when 16#18e6# => read_data_o <= x"0000";
				when 16#18e7# => read_data_o <= x"0000";
				when 16#18e8# => read_data_o <= x"0000";
				when 16#18e9# => read_data_o <= x"0000";
				when 16#18ea# => read_data_o <= x"0000";
				when 16#18eb# => read_data_o <= x"0000";
				when 16#18ec# => read_data_o <= x"0000";
				when 16#18ed# => read_data_o <= x"0000";
				when 16#18ee# => read_data_o <= x"0000";
				when 16#18ef# => read_data_o <= x"0000";
				when 16#18f0# => read_data_o <= x"0000";
				when 16#18f1# => read_data_o <= x"0000";
				when 16#18f2# => read_data_o <= x"0000";
				when 16#18f3# => read_data_o <= x"0000";
				when 16#18f4# => read_data_o <= x"0000";
				when 16#18f5# => read_data_o <= x"0000";
				when 16#18f6# => read_data_o <= x"0000";
				when 16#18f7# => read_data_o <= x"0000";
				when 16#18f8# => read_data_o <= x"0000";
				when 16#18f9# => read_data_o <= x"0000";
				when 16#18fa# => read_data_o <= x"0000";
				when 16#18fb# => read_data_o <= x"0000";
				when 16#18fc# => read_data_o <= x"0000";
				when 16#18fd# => read_data_o <= x"0000";
				when 16#18fe# => read_data_o <= x"0000";
				when 16#18ff# => read_data_o <= x"0000";
				when 16#1900# => read_data_o <= x"0000";
				when 16#1901# => read_data_o <= x"0000";
				when 16#1902# => read_data_o <= x"0000";
				when 16#1903# => read_data_o <= x"0000";
				when 16#1904# => read_data_o <= x"0000";
				when 16#1905# => read_data_o <= x"0000";
				when 16#1906# => read_data_o <= x"0000";
				when 16#1907# => read_data_o <= x"0000";
				when 16#1908# => read_data_o <= x"0000";
				when 16#1909# => read_data_o <= x"0000";
				when 16#190a# => read_data_o <= x"0000";
				when 16#190b# => read_data_o <= x"0000";
				when 16#190c# => read_data_o <= x"0000";
				when 16#190d# => read_data_o <= x"0000";
				when 16#190e# => read_data_o <= x"0000";
				when 16#190f# => read_data_o <= x"0000";
				when 16#1910# => read_data_o <= x"0000";
				when 16#1911# => read_data_o <= x"0000";
				when 16#1912# => read_data_o <= x"0000";
				when 16#1913# => read_data_o <= x"0000";
				when 16#1914# => read_data_o <= x"0000";
				when 16#1915# => read_data_o <= x"0000";
				when 16#1916# => read_data_o <= x"0000";
				when 16#1917# => read_data_o <= x"0000";
				when 16#1918# => read_data_o <= x"0000";
				when 16#1919# => read_data_o <= x"0000";
				when 16#191a# => read_data_o <= x"0000";
				when 16#191b# => read_data_o <= x"0000";
				when 16#191c# => read_data_o <= x"0000";
				when 16#191d# => read_data_o <= x"0000";
				when 16#191e# => read_data_o <= x"0000";
				when 16#191f# => read_data_o <= x"0000";
				when 16#1920# => read_data_o <= x"0000";
				when 16#1921# => read_data_o <= x"0000";
				when 16#1922# => read_data_o <= x"0000";
				when 16#1923# => read_data_o <= x"0000";
				when 16#1924# => read_data_o <= x"0000";
				when 16#1925# => read_data_o <= x"0000";
				when 16#1926# => read_data_o <= x"0000";
				when 16#1927# => read_data_o <= x"0000";
				when 16#1928# => read_data_o <= x"0000";
				when 16#1929# => read_data_o <= x"0000";
				when 16#192a# => read_data_o <= x"0000";
				when 16#192b# => read_data_o <= x"0000";
				when 16#192c# => read_data_o <= x"0000";
				when 16#192d# => read_data_o <= x"0000";
				when 16#192e# => read_data_o <= x"0000";
				when 16#192f# => read_data_o <= x"0000";
				when 16#1930# => read_data_o <= x"0000";
				when 16#1931# => read_data_o <= x"0000";
				when 16#1932# => read_data_o <= x"0000";
				when 16#1933# => read_data_o <= x"0000";
				when 16#1934# => read_data_o <= x"0000";
				when 16#1935# => read_data_o <= x"0000";
				when 16#1936# => read_data_o <= x"0000";
				when 16#1937# => read_data_o <= x"0000";
				when 16#1938# => read_data_o <= x"0000";
				when 16#1939# => read_data_o <= x"0000";
				when 16#193a# => read_data_o <= x"0000";
				when 16#193b# => read_data_o <= x"0000";
				when 16#193c# => read_data_o <= x"0000";
				when 16#193d# => read_data_o <= x"0000";
				when 16#193e# => read_data_o <= x"0000";
				when 16#193f# => read_data_o <= x"0000";
				when 16#1940# => read_data_o <= x"0000";
				when 16#1941# => read_data_o <= x"0000";
				when 16#1942# => read_data_o <= x"0000";
				when 16#1943# => read_data_o <= x"0000";
				when 16#1944# => read_data_o <= x"0000";
				when 16#1945# => read_data_o <= x"0000";
				when 16#1946# => read_data_o <= x"0000";
				when 16#1947# => read_data_o <= x"0000";
				when 16#1948# => read_data_o <= x"0000";
				when 16#1949# => read_data_o <= x"0000";
				when 16#194a# => read_data_o <= x"0000";
				when 16#194b# => read_data_o <= x"0000";
				when 16#194c# => read_data_o <= x"0000";
				when 16#194d# => read_data_o <= x"0000";
				when 16#194e# => read_data_o <= x"0000";
				when 16#194f# => read_data_o <= x"0000";
				when 16#1950# => read_data_o <= x"0000";
				when 16#1951# => read_data_o <= x"0000";
				when 16#1952# => read_data_o <= x"0000";
				when 16#1953# => read_data_o <= x"0000";
				when 16#1954# => read_data_o <= x"0000";
				when 16#1955# => read_data_o <= x"0000";
				when 16#1956# => read_data_o <= x"0000";
				when 16#1957# => read_data_o <= x"0000";
				when 16#1958# => read_data_o <= x"0000";
				when 16#1959# => read_data_o <= x"0000";
				when 16#195a# => read_data_o <= x"0000";
				when 16#195b# => read_data_o <= x"0000";
				when 16#195c# => read_data_o <= x"0000";
				when 16#195d# => read_data_o <= x"0000";
				when 16#195e# => read_data_o <= x"0000";
				when 16#195f# => read_data_o <= x"0000";
				when 16#1960# => read_data_o <= x"0000";
				when 16#1961# => read_data_o <= x"0000";
				when 16#1962# => read_data_o <= x"0000";
				when 16#1963# => read_data_o <= x"0000";
				when 16#1964# => read_data_o <= x"0000";
				when 16#1965# => read_data_o <= x"0000";
				when 16#1966# => read_data_o <= x"0000";
				when 16#1967# => read_data_o <= x"0000";
				when 16#1968# => read_data_o <= x"0000";
				when 16#1969# => read_data_o <= x"0000";
				when 16#196a# => read_data_o <= x"0000";
				when 16#196b# => read_data_o <= x"0000";
				when 16#196c# => read_data_o <= x"0000";
				when 16#196d# => read_data_o <= x"0000";
				when 16#196e# => read_data_o <= x"0000";
				when 16#196f# => read_data_o <= x"0000";
				when 16#1970# => read_data_o <= x"0000";
				when 16#1971# => read_data_o <= x"0000";
				when 16#1972# => read_data_o <= x"0000";
				when 16#1973# => read_data_o <= x"0000";
				when 16#1974# => read_data_o <= x"0000";
				when 16#1975# => read_data_o <= x"0000";
				when 16#1976# => read_data_o <= x"0000";
				when 16#1977# => read_data_o <= x"0000";
				when 16#1978# => read_data_o <= x"0000";
				when 16#1979# => read_data_o <= x"0000";
				when 16#197a# => read_data_o <= x"0000";
				when 16#197b# => read_data_o <= x"0000";
				when 16#197c# => read_data_o <= x"0000";
				when 16#197d# => read_data_o <= x"0000";
				when 16#197e# => read_data_o <= x"0000";
				when 16#197f# => read_data_o <= x"0000";
				when 16#1980# => read_data_o <= x"0000";
				when 16#1981# => read_data_o <= x"0000";
				when 16#1982# => read_data_o <= x"0000";
				when 16#1983# => read_data_o <= x"0000";
				when 16#1984# => read_data_o <= x"0000";
				when 16#1985# => read_data_o <= x"0000";
				when 16#1986# => read_data_o <= x"0000";
				when 16#1987# => read_data_o <= x"0000";
				when 16#1988# => read_data_o <= x"0000";
				when 16#1989# => read_data_o <= x"0000";
				when 16#198a# => read_data_o <= x"0000";
				when 16#198b# => read_data_o <= x"0000";
				when 16#198c# => read_data_o <= x"0000";
				when 16#198d# => read_data_o <= x"0000";
				when 16#198e# => read_data_o <= x"0000";
				when 16#198f# => read_data_o <= x"0000";
				when 16#1990# => read_data_o <= x"0000";
				when 16#1991# => read_data_o <= x"0000";
				when 16#1992# => read_data_o <= x"0000";
				when 16#1993# => read_data_o <= x"0000";
				when 16#1994# => read_data_o <= x"0000";
				when 16#1995# => read_data_o <= x"0000";
				when 16#1996# => read_data_o <= x"0000";
				when 16#1997# => read_data_o <= x"0000";
				when 16#1998# => read_data_o <= x"0000";
				when 16#1999# => read_data_o <= x"0000";
				when 16#199a# => read_data_o <= x"0000";
				when 16#199b# => read_data_o <= x"0000";
				when 16#199c# => read_data_o <= x"0000";
				when 16#199d# => read_data_o <= x"0000";
				when 16#199e# => read_data_o <= x"0000";
				when 16#199f# => read_data_o <= x"0000";
				when 16#19a0# => read_data_o <= x"0000";
				when 16#19a1# => read_data_o <= x"0000";
				when 16#19a2# => read_data_o <= x"0000";
				when 16#19a3# => read_data_o <= x"0000";
				when 16#19a4# => read_data_o <= x"0000";
				when 16#19a5# => read_data_o <= x"0000";
				when 16#19a6# => read_data_o <= x"0000";
				when 16#19a7# => read_data_o <= x"0000";
				when 16#19a8# => read_data_o <= x"0000";
				when 16#19a9# => read_data_o <= x"0000";
				when 16#19aa# => read_data_o <= x"0000";
				when 16#19ab# => read_data_o <= x"0000";
				when 16#19ac# => read_data_o <= x"0000";
				when 16#19ad# => read_data_o <= x"0000";
				when 16#19ae# => read_data_o <= x"0000";
				when 16#19af# => read_data_o <= x"0000";
				when 16#19b0# => read_data_o <= x"0000";
				when 16#19b1# => read_data_o <= x"0000";
				when 16#19b2# => read_data_o <= x"0000";
				when 16#19b3# => read_data_o <= x"0000";
				when 16#19b4# => read_data_o <= x"0000";
				when 16#19b5# => read_data_o <= x"0000";
				when 16#19b6# => read_data_o <= x"0000";
				when 16#19b7# => read_data_o <= x"0000";
				when 16#19b8# => read_data_o <= x"0000";
				when 16#19b9# => read_data_o <= x"0000";
				when 16#19ba# => read_data_o <= x"0000";
				when 16#19bb# => read_data_o <= x"0000";
				when 16#19bc# => read_data_o <= x"0000";
				when 16#19bd# => read_data_o <= x"0000";
				when 16#19be# => read_data_o <= x"0000";
				when 16#19bf# => read_data_o <= x"0000";
				when 16#19c0# => read_data_o <= x"0000";
				when 16#19c1# => read_data_o <= x"0000";
				when 16#19c2# => read_data_o <= x"0000";
				when 16#19c3# => read_data_o <= x"0000";
				when 16#19c4# => read_data_o <= x"0000";
				when 16#19c5# => read_data_o <= x"0000";
				when 16#19c6# => read_data_o <= x"0000";
				when 16#19c7# => read_data_o <= x"0000";
				when 16#19c8# => read_data_o <= x"0000";
				when 16#19c9# => read_data_o <= x"0000";
				when 16#19ca# => read_data_o <= x"0000";
				when 16#19cb# => read_data_o <= x"0000";
				when 16#19cc# => read_data_o <= x"0000";
				when 16#19cd# => read_data_o <= x"0000";
				when 16#19ce# => read_data_o <= x"0000";
				when 16#19cf# => read_data_o <= x"0000";
				when 16#19d0# => read_data_o <= x"0000";
				when 16#19d1# => read_data_o <= x"0000";
				when 16#19d2# => read_data_o <= x"0000";
				when 16#19d3# => read_data_o <= x"0000";
				when 16#19d4# => read_data_o <= x"0000";
				when 16#19d5# => read_data_o <= x"0000";
				when 16#19d6# => read_data_o <= x"0000";
				when 16#19d7# => read_data_o <= x"0000";
				when 16#19d8# => read_data_o <= x"0000";
				when 16#19d9# => read_data_o <= x"0000";
				when 16#19da# => read_data_o <= x"0000";
				when 16#19db# => read_data_o <= x"0000";
				when 16#19dc# => read_data_o <= x"0000";
				when 16#19dd# => read_data_o <= x"0000";
				when 16#19de# => read_data_o <= x"0000";
				when 16#19df# => read_data_o <= x"0000";
				when 16#19e0# => read_data_o <= x"0000";
				when 16#19e1# => read_data_o <= x"0000";
				when 16#19e2# => read_data_o <= x"0000";
				when 16#19e3# => read_data_o <= x"0000";
				when 16#19e4# => read_data_o <= x"0000";
				when 16#19e5# => read_data_o <= x"0000";
				when 16#19e6# => read_data_o <= x"0000";
				when 16#19e7# => read_data_o <= x"0000";
				when 16#19e8# => read_data_o <= x"0000";
				when 16#19e9# => read_data_o <= x"0000";
				when 16#19ea# => read_data_o <= x"0000";
				when 16#19eb# => read_data_o <= x"0000";
				when 16#19ec# => read_data_o <= x"0000";
				when 16#19ed# => read_data_o <= x"0000";
				when 16#19ee# => read_data_o <= x"0000";
				when 16#19ef# => read_data_o <= x"0000";
				when 16#19f0# => read_data_o <= x"0000";
				when 16#19f1# => read_data_o <= x"0000";
				when 16#19f2# => read_data_o <= x"0000";
				when 16#19f3# => read_data_o <= x"0000";
				when 16#19f4# => read_data_o <= x"0000";
				when 16#19f5# => read_data_o <= x"0000";
				when 16#19f6# => read_data_o <= x"0000";
				when 16#19f7# => read_data_o <= x"0000";
				when 16#19f8# => read_data_o <= x"0000";
				when 16#19f9# => read_data_o <= x"0000";
				when 16#19fa# => read_data_o <= x"0000";
				when 16#19fb# => read_data_o <= x"0000";
				when 16#19fc# => read_data_o <= x"0000";
				when 16#19fd# => read_data_o <= x"0000";
				when 16#19fe# => read_data_o <= x"0000";
				when 16#19ff# => read_data_o <= x"0000";
				when 16#1a00# => read_data_o <= x"0000";
				when 16#1a01# => read_data_o <= x"0000";
				when 16#1a02# => read_data_o <= x"0000";
				when 16#1a03# => read_data_o <= x"0000";
				when 16#1a04# => read_data_o <= x"0000";
				when 16#1a05# => read_data_o <= x"0000";
				when 16#1a06# => read_data_o <= x"0000";
				when 16#1a07# => read_data_o <= x"0000";
				when 16#1a08# => read_data_o <= x"0000";
				when 16#1a09# => read_data_o <= x"0000";
				when 16#1a0a# => read_data_o <= x"0000";
				when 16#1a0b# => read_data_o <= x"0000";
				when 16#1a0c# => read_data_o <= x"0000";
				when 16#1a0d# => read_data_o <= x"0000";
				when 16#1a0e# => read_data_o <= x"0000";
				when 16#1a0f# => read_data_o <= x"0000";
				when 16#1a10# => read_data_o <= x"0000";
				when 16#1a11# => read_data_o <= x"0000";
				when 16#1a12# => read_data_o <= x"0000";
				when 16#1a13# => read_data_o <= x"0000";
				when 16#1a14# => read_data_o <= x"0000";
				when 16#1a15# => read_data_o <= x"0000";
				when 16#1a16# => read_data_o <= x"0000";
				when 16#1a17# => read_data_o <= x"0000";
				when 16#1a18# => read_data_o <= x"0000";
				when 16#1a19# => read_data_o <= x"0000";
				when 16#1a1a# => read_data_o <= x"0000";
				when 16#1a1b# => read_data_o <= x"0000";
				when 16#1a1c# => read_data_o <= x"0000";
				when 16#1a1d# => read_data_o <= x"0000";
				when 16#1a1e# => read_data_o <= x"0000";
				when 16#1a1f# => read_data_o <= x"0000";
				when 16#1a20# => read_data_o <= x"0000";
				when 16#1a21# => read_data_o <= x"0000";
				when 16#1a22# => read_data_o <= x"0000";
				when 16#1a23# => read_data_o <= x"0000";
				when 16#1a24# => read_data_o <= x"0000";
				when 16#1a25# => read_data_o <= x"0000";
				when 16#1a26# => read_data_o <= x"0000";
				when 16#1a27# => read_data_o <= x"0000";
				when 16#1a28# => read_data_o <= x"0000";
				when 16#1a29# => read_data_o <= x"0000";
				when 16#1a2a# => read_data_o <= x"0000";
				when 16#1a2b# => read_data_o <= x"0000";
				when 16#1a2c# => read_data_o <= x"0000";
				when 16#1a2d# => read_data_o <= x"0000";
				when 16#1a2e# => read_data_o <= x"0000";
				when 16#1a2f# => read_data_o <= x"0000";
				when 16#1a30# => read_data_o <= x"0000";
				when 16#1a31# => read_data_o <= x"0000";
				when 16#1a32# => read_data_o <= x"0000";
				when 16#1a33# => read_data_o <= x"0000";
				when 16#1a34# => read_data_o <= x"0000";
				when 16#1a35# => read_data_o <= x"0000";
				when 16#1a36# => read_data_o <= x"0000";
				when 16#1a37# => read_data_o <= x"0000";
				when 16#1a38# => read_data_o <= x"0000";
				when 16#1a39# => read_data_o <= x"0000";
				when 16#1a3a# => read_data_o <= x"0000";
				when 16#1a3b# => read_data_o <= x"0000";
				when 16#1a3c# => read_data_o <= x"0000";
				when 16#1a3d# => read_data_o <= x"0000";
				when 16#1a3e# => read_data_o <= x"0000";
				when 16#1a3f# => read_data_o <= x"0000";
				when 16#1a40# => read_data_o <= x"0000";
				when 16#1a41# => read_data_o <= x"0000";
				when 16#1a42# => read_data_o <= x"0000";
				when 16#1a43# => read_data_o <= x"0000";
				when 16#1a44# => read_data_o <= x"0000";
				when 16#1a45# => read_data_o <= x"0000";
				when 16#1a46# => read_data_o <= x"0000";
				when 16#1a47# => read_data_o <= x"0000";
				when 16#1a48# => read_data_o <= x"0000";
				when 16#1a49# => read_data_o <= x"0000";
				when 16#1a4a# => read_data_o <= x"0000";
				when 16#1a4b# => read_data_o <= x"0000";
				when 16#1a4c# => read_data_o <= x"0000";
				when 16#1a4d# => read_data_o <= x"0000";
				when 16#1a4e# => read_data_o <= x"0000";
				when 16#1a4f# => read_data_o <= x"0000";
				when 16#1a50# => read_data_o <= x"0000";
				when 16#1a51# => read_data_o <= x"0000";
				when 16#1a52# => read_data_o <= x"0000";
				when 16#1a53# => read_data_o <= x"0000";
				when 16#1a54# => read_data_o <= x"0000";
				when 16#1a55# => read_data_o <= x"0000";
				when 16#1a56# => read_data_o <= x"0000";
				when 16#1a57# => read_data_o <= x"0000";
				when 16#1a58# => read_data_o <= x"0000";
				when 16#1a59# => read_data_o <= x"0000";
				when 16#1a5a# => read_data_o <= x"0000";
				when 16#1a5b# => read_data_o <= x"0000";
				when 16#1a5c# => read_data_o <= x"0000";
				when 16#1a5d# => read_data_o <= x"0000";
				when 16#1a5e# => read_data_o <= x"0000";
				when 16#1a5f# => read_data_o <= x"0000";
				when 16#1a60# => read_data_o <= x"0000";
				when 16#1a61# => read_data_o <= x"0000";
				when 16#1a62# => read_data_o <= x"0000";
				when 16#1a63# => read_data_o <= x"0000";
				when 16#1a64# => read_data_o <= x"0000";
				when 16#1a65# => read_data_o <= x"0000";
				when 16#1a66# => read_data_o <= x"0000";
				when 16#1a67# => read_data_o <= x"0000";
				when 16#1a68# => read_data_o <= x"0000";
				when 16#1a69# => read_data_o <= x"0000";
				when 16#1a6a# => read_data_o <= x"0000";
				when 16#1a6b# => read_data_o <= x"0000";
				when 16#1a6c# => read_data_o <= x"0000";
				when 16#1a6d# => read_data_o <= x"0000";
				when 16#1a6e# => read_data_o <= x"0000";
				when 16#1a6f# => read_data_o <= x"0000";
				when 16#1a70# => read_data_o <= x"0000";
				when 16#1a71# => read_data_o <= x"0000";
				when 16#1a72# => read_data_o <= x"0000";
				when 16#1a73# => read_data_o <= x"0000";
				when 16#1a74# => read_data_o <= x"0000";
				when 16#1a75# => read_data_o <= x"0000";
				when 16#1a76# => read_data_o <= x"0000";
				when 16#1a77# => read_data_o <= x"0000";
				when 16#1a78# => read_data_o <= x"0000";
				when 16#1a79# => read_data_o <= x"0000";
				when 16#1a7a# => read_data_o <= x"0000";
				when 16#1a7b# => read_data_o <= x"0000";
				when 16#1a7c# => read_data_o <= x"0000";
				when 16#1a7d# => read_data_o <= x"0000";
				when 16#1a7e# => read_data_o <= x"0000";
				when 16#1a7f# => read_data_o <= x"0000";
				when 16#1a80# => read_data_o <= x"0000";
				when 16#1a81# => read_data_o <= x"0000";
				when 16#1a82# => read_data_o <= x"0000";
				when 16#1a83# => read_data_o <= x"0000";
				when 16#1a84# => read_data_o <= x"0000";
				when 16#1a85# => read_data_o <= x"0000";
				when 16#1a86# => read_data_o <= x"0000";
				when 16#1a87# => read_data_o <= x"0000";
				when 16#1a88# => read_data_o <= x"0000";
				when 16#1a89# => read_data_o <= x"0000";
				when 16#1a8a# => read_data_o <= x"0000";
				when 16#1a8b# => read_data_o <= x"0000";
				when 16#1a8c# => read_data_o <= x"0000";
				when 16#1a8d# => read_data_o <= x"0000";
				when 16#1a8e# => read_data_o <= x"0000";
				when 16#1a8f# => read_data_o <= x"0000";
				when 16#1a90# => read_data_o <= x"0000";
				when 16#1a91# => read_data_o <= x"0000";
				when 16#1a92# => read_data_o <= x"0000";
				when 16#1a93# => read_data_o <= x"0000";
				when 16#1a94# => read_data_o <= x"0000";
				when 16#1a95# => read_data_o <= x"0000";
				when 16#1a96# => read_data_o <= x"0000";
				when 16#1a97# => read_data_o <= x"0000";
				when 16#1a98# => read_data_o <= x"0000";
				when 16#1a99# => read_data_o <= x"0000";
				when 16#1a9a# => read_data_o <= x"0000";
				when 16#1a9b# => read_data_o <= x"0000";
				when 16#1a9c# => read_data_o <= x"0000";
				when 16#1a9d# => read_data_o <= x"0000";
				when 16#1a9e# => read_data_o <= x"0000";
				when 16#1a9f# => read_data_o <= x"0000";
				when 16#1aa0# => read_data_o <= x"0000";
				when 16#1aa1# => read_data_o <= x"0000";
				when 16#1aa2# => read_data_o <= x"0000";
				when 16#1aa3# => read_data_o <= x"0000";
				when 16#1aa4# => read_data_o <= x"0000";
				when 16#1aa5# => read_data_o <= x"0000";
				when 16#1aa6# => read_data_o <= x"0000";
				when 16#1aa7# => read_data_o <= x"0000";
				when 16#1aa8# => read_data_o <= x"0000";
				when 16#1aa9# => read_data_o <= x"0000";
				when 16#1aaa# => read_data_o <= x"0000";
				when 16#1aab# => read_data_o <= x"0000";
				when 16#1aac# => read_data_o <= x"0000";
				when 16#1aad# => read_data_o <= x"0000";
				when 16#1aae# => read_data_o <= x"0000";
				when 16#1aaf# => read_data_o <= x"0000";
				when 16#1ab0# => read_data_o <= x"0000";
				when 16#1ab1# => read_data_o <= x"0000";
				when 16#1ab2# => read_data_o <= x"0000";
				when 16#1ab3# => read_data_o <= x"0000";
				when 16#1ab4# => read_data_o <= x"0000";
				when 16#1ab5# => read_data_o <= x"0000";
				when 16#1ab6# => read_data_o <= x"0000";
				when 16#1ab7# => read_data_o <= x"0000";
				when 16#1ab8# => read_data_o <= x"0000";
				when 16#1ab9# => read_data_o <= x"0000";
				when 16#1aba# => read_data_o <= x"0000";
				when 16#1abb# => read_data_o <= x"0000";
				when 16#1abc# => read_data_o <= x"0000";
				when 16#1abd# => read_data_o <= x"0000";
				when 16#1abe# => read_data_o <= x"0000";
				when 16#1abf# => read_data_o <= x"0000";
				when 16#1ac0# => read_data_o <= x"0000";
				when 16#1ac1# => read_data_o <= x"0000";
				when 16#1ac2# => read_data_o <= x"0000";
				when 16#1ac3# => read_data_o <= x"0000";
				when 16#1ac4# => read_data_o <= x"0000";
				when 16#1ac5# => read_data_o <= x"0000";
				when 16#1ac6# => read_data_o <= x"0000";
				when 16#1ac7# => read_data_o <= x"0000";
				when 16#1ac8# => read_data_o <= x"0000";
				when 16#1ac9# => read_data_o <= x"0000";
				when 16#1aca# => read_data_o <= x"0000";
				when 16#1acb# => read_data_o <= x"0000";
				when 16#1acc# => read_data_o <= x"0000";
				when 16#1acd# => read_data_o <= x"0000";
				when 16#1ace# => read_data_o <= x"0000";
				when 16#1acf# => read_data_o <= x"0000";
				when 16#1ad0# => read_data_o <= x"0000";
				when 16#1ad1# => read_data_o <= x"0000";
				when 16#1ad2# => read_data_o <= x"0000";
				when 16#1ad3# => read_data_o <= x"0000";
				when 16#1ad4# => read_data_o <= x"0000";
				when 16#1ad5# => read_data_o <= x"0000";
				when 16#1ad6# => read_data_o <= x"0000";
				when 16#1ad7# => read_data_o <= x"0000";
				when 16#1ad8# => read_data_o <= x"0000";
				when 16#1ad9# => read_data_o <= x"0000";
				when 16#1ada# => read_data_o <= x"0000";
				when 16#1adb# => read_data_o <= x"0000";
				when 16#1adc# => read_data_o <= x"0000";
				when 16#1add# => read_data_o <= x"0000";
				when 16#1ade# => read_data_o <= x"0000";
				when 16#1adf# => read_data_o <= x"0000";
				when 16#1ae0# => read_data_o <= x"0000";
				when 16#1ae1# => read_data_o <= x"0000";
				when 16#1ae2# => read_data_o <= x"0000";
				when 16#1ae3# => read_data_o <= x"0000";
				when 16#1ae4# => read_data_o <= x"0000";
				when 16#1ae5# => read_data_o <= x"0000";
				when 16#1ae6# => read_data_o <= x"0000";
				when 16#1ae7# => read_data_o <= x"0000";
				when 16#1ae8# => read_data_o <= x"0000";
				when 16#1ae9# => read_data_o <= x"0000";
				when 16#1aea# => read_data_o <= x"0000";
				when 16#1aeb# => read_data_o <= x"0000";
				when 16#1aec# => read_data_o <= x"0000";
				when 16#1aed# => read_data_o <= x"0000";
				when 16#1aee# => read_data_o <= x"0000";
				when 16#1aef# => read_data_o <= x"0000";
				when 16#1af0# => read_data_o <= x"0000";
				when 16#1af1# => read_data_o <= x"0000";
				when 16#1af2# => read_data_o <= x"0000";
				when 16#1af3# => read_data_o <= x"0000";
				when 16#1af4# => read_data_o <= x"0000";
				when 16#1af5# => read_data_o <= x"0000";
				when 16#1af6# => read_data_o <= x"0000";
				when 16#1af7# => read_data_o <= x"0000";
				when 16#1af8# => read_data_o <= x"0000";
				when 16#1af9# => read_data_o <= x"0000";
				when 16#1afa# => read_data_o <= x"0000";
				when 16#1afb# => read_data_o <= x"0000";
				when 16#1afc# => read_data_o <= x"0000";
				when 16#1afd# => read_data_o <= x"0000";
				when 16#1afe# => read_data_o <= x"0000";
				when 16#1aff# => read_data_o <= x"0000";
				when 16#1b00# => read_data_o <= x"0000";
				when 16#1b01# => read_data_o <= x"0000";
				when 16#1b02# => read_data_o <= x"0000";
				when 16#1b03# => read_data_o <= x"0000";
				when 16#1b04# => read_data_o <= x"0000";
				when 16#1b05# => read_data_o <= x"0000";
				when 16#1b06# => read_data_o <= x"0000";
				when 16#1b07# => read_data_o <= x"0000";
				when 16#1b08# => read_data_o <= x"0000";
				when 16#1b09# => read_data_o <= x"0000";
				when 16#1b0a# => read_data_o <= x"0000";
				when 16#1b0b# => read_data_o <= x"0000";
				when 16#1b0c# => read_data_o <= x"0000";
				when 16#1b0d# => read_data_o <= x"0000";
				when 16#1b0e# => read_data_o <= x"0000";
				when 16#1b0f# => read_data_o <= x"0000";
				when 16#1b10# => read_data_o <= x"0000";
				when 16#1b11# => read_data_o <= x"0000";
				when 16#1b12# => read_data_o <= x"0000";
				when 16#1b13# => read_data_o <= x"0000";
				when 16#1b14# => read_data_o <= x"0000";
				when 16#1b15# => read_data_o <= x"0000";
				when 16#1b16# => read_data_o <= x"0000";
				when 16#1b17# => read_data_o <= x"0000";
				when 16#1b18# => read_data_o <= x"0000";
				when 16#1b19# => read_data_o <= x"0000";
				when 16#1b1a# => read_data_o <= x"0000";
				when 16#1b1b# => read_data_o <= x"0000";
				when 16#1b1c# => read_data_o <= x"0000";
				when 16#1b1d# => read_data_o <= x"0000";
				when 16#1b1e# => read_data_o <= x"0000";
				when 16#1b1f# => read_data_o <= x"0000";
				when 16#1b20# => read_data_o <= x"0000";
				when 16#1b21# => read_data_o <= x"0000";
				when 16#1b22# => read_data_o <= x"0000";
				when 16#1b23# => read_data_o <= x"0000";
				when 16#1b24# => read_data_o <= x"0000";
				when 16#1b25# => read_data_o <= x"0000";
				when 16#1b26# => read_data_o <= x"0000";
				when 16#1b27# => read_data_o <= x"0000";
				when 16#1b28# => read_data_o <= x"0000";
				when 16#1b29# => read_data_o <= x"0000";
				when 16#1b2a# => read_data_o <= x"0000";
				when 16#1b2b# => read_data_o <= x"0000";
				when 16#1b2c# => read_data_o <= x"0000";
				when 16#1b2d# => read_data_o <= x"0000";
				when 16#1b2e# => read_data_o <= x"0000";
				when 16#1b2f# => read_data_o <= x"0000";
				when 16#1b30# => read_data_o <= x"0000";
				when 16#1b31# => read_data_o <= x"0000";
				when 16#1b32# => read_data_o <= x"0000";
				when 16#1b33# => read_data_o <= x"0000";
				when 16#1b34# => read_data_o <= x"0000";
				when 16#1b35# => read_data_o <= x"0000";
				when 16#1b36# => read_data_o <= x"0000";
				when 16#1b37# => read_data_o <= x"0000";
				when 16#1b38# => read_data_o <= x"0000";
				when 16#1b39# => read_data_o <= x"0000";
				when 16#1b3a# => read_data_o <= x"0000";
				when 16#1b3b# => read_data_o <= x"0000";
				when 16#1b3c# => read_data_o <= x"0000";
				when 16#1b3d# => read_data_o <= x"0000";
				when 16#1b3e# => read_data_o <= x"0000";
				when 16#1b3f# => read_data_o <= x"0000";
				when 16#1b40# => read_data_o <= x"0000";
				when 16#1b41# => read_data_o <= x"0000";
				when 16#1b42# => read_data_o <= x"0000";
				when 16#1b43# => read_data_o <= x"0000";
				when 16#1b44# => read_data_o <= x"0000";
				when 16#1b45# => read_data_o <= x"0000";
				when 16#1b46# => read_data_o <= x"0000";
				when 16#1b47# => read_data_o <= x"0000";
				when 16#1b48# => read_data_o <= x"0000";
				when 16#1b49# => read_data_o <= x"0000";
				when 16#1b4a# => read_data_o <= x"0000";
				when 16#1b4b# => read_data_o <= x"0000";
				when 16#1b4c# => read_data_o <= x"0000";
				when 16#1b4d# => read_data_o <= x"0000";
				when 16#1b4e# => read_data_o <= x"0000";
				when 16#1b4f# => read_data_o <= x"0000";
				when 16#1b50# => read_data_o <= x"0000";
				when 16#1b51# => read_data_o <= x"0000";
				when 16#1b52# => read_data_o <= x"0000";
				when 16#1b53# => read_data_o <= x"0000";
				when 16#1b54# => read_data_o <= x"0000";
				when 16#1b55# => read_data_o <= x"0000";
				when 16#1b56# => read_data_o <= x"0000";
				when 16#1b57# => read_data_o <= x"0000";
				when 16#1b58# => read_data_o <= x"0000";
				when 16#1b59# => read_data_o <= x"0000";
				when 16#1b5a# => read_data_o <= x"0000";
				when 16#1b5b# => read_data_o <= x"0000";
				when 16#1b5c# => read_data_o <= x"0000";
				when 16#1b5d# => read_data_o <= x"0000";
				when 16#1b5e# => read_data_o <= x"0000";
				when 16#1b5f# => read_data_o <= x"0000";
				when 16#1b60# => read_data_o <= x"0000";
				when 16#1b61# => read_data_o <= x"0000";
				when 16#1b62# => read_data_o <= x"0000";
				when 16#1b63# => read_data_o <= x"0000";
				when 16#1b64# => read_data_o <= x"0000";
				when 16#1b65# => read_data_o <= x"0000";
				when 16#1b66# => read_data_o <= x"0000";
				when 16#1b67# => read_data_o <= x"0000";
				when 16#1b68# => read_data_o <= x"0000";
				when 16#1b69# => read_data_o <= x"0000";
				when 16#1b6a# => read_data_o <= x"0000";
				when 16#1b6b# => read_data_o <= x"0000";
				when 16#1b6c# => read_data_o <= x"0000";
				when 16#1b6d# => read_data_o <= x"0000";
				when 16#1b6e# => read_data_o <= x"0000";
				when 16#1b6f# => read_data_o <= x"0000";
				when 16#1b70# => read_data_o <= x"0000";
				when 16#1b71# => read_data_o <= x"0000";
				when 16#1b72# => read_data_o <= x"0000";
				when 16#1b73# => read_data_o <= x"0000";
				when 16#1b74# => read_data_o <= x"0000";
				when 16#1b75# => read_data_o <= x"0000";
				when 16#1b76# => read_data_o <= x"0000";
				when 16#1b77# => read_data_o <= x"0000";
				when 16#1b78# => read_data_o <= x"0000";
				when 16#1b79# => read_data_o <= x"0000";
				when 16#1b7a# => read_data_o <= x"0000";
				when 16#1b7b# => read_data_o <= x"0000";
				when 16#1b7c# => read_data_o <= x"0000";
				when 16#1b7d# => read_data_o <= x"0000";
				when 16#1b7e# => read_data_o <= x"0000";
				when 16#1b7f# => read_data_o <= x"0000";
				when 16#1b80# => read_data_o <= x"0000";
				when 16#1b81# => read_data_o <= x"0000";
				when 16#1b82# => read_data_o <= x"0000";
				when 16#1b83# => read_data_o <= x"0000";
				when 16#1b84# => read_data_o <= x"0000";
				when 16#1b85# => read_data_o <= x"0000";
				when 16#1b86# => read_data_o <= x"0000";
				when 16#1b87# => read_data_o <= x"0000";
				when 16#1b88# => read_data_o <= x"0000";
				when 16#1b89# => read_data_o <= x"0000";
				when 16#1b8a# => read_data_o <= x"0000";
				when 16#1b8b# => read_data_o <= x"0000";
				when 16#1b8c# => read_data_o <= x"0000";
				when 16#1b8d# => read_data_o <= x"0000";
				when 16#1b8e# => read_data_o <= x"0000";
				when 16#1b8f# => read_data_o <= x"0000";
				when 16#1b90# => read_data_o <= x"0000";
				when 16#1b91# => read_data_o <= x"0000";
				when 16#1b92# => read_data_o <= x"0000";
				when 16#1b93# => read_data_o <= x"0000";
				when 16#1b94# => read_data_o <= x"0000";
				when 16#1b95# => read_data_o <= x"0000";
				when 16#1b96# => read_data_o <= x"0000";
				when 16#1b97# => read_data_o <= x"0000";
				when 16#1b98# => read_data_o <= x"0000";
				when 16#1b99# => read_data_o <= x"0000";
				when 16#1b9a# => read_data_o <= x"0000";
				when 16#1b9b# => read_data_o <= x"0000";
				when 16#1b9c# => read_data_o <= x"0000";
				when 16#1b9d# => read_data_o <= x"0000";
				when 16#1b9e# => read_data_o <= x"0000";
				when 16#1b9f# => read_data_o <= x"0000";
				when 16#1ba0# => read_data_o <= x"0000";
				when 16#1ba1# => read_data_o <= x"0000";
				when 16#1ba2# => read_data_o <= x"0000";
				when 16#1ba3# => read_data_o <= x"0000";
				when 16#1ba4# => read_data_o <= x"0000";
				when 16#1ba5# => read_data_o <= x"0000";
				when 16#1ba6# => read_data_o <= x"0000";
				when 16#1ba7# => read_data_o <= x"0000";
				when 16#1ba8# => read_data_o <= x"0000";
				when 16#1ba9# => read_data_o <= x"0000";
				when 16#1baa# => read_data_o <= x"0000";
				when 16#1bab# => read_data_o <= x"0000";
				when 16#1bac# => read_data_o <= x"0000";
				when 16#1bad# => read_data_o <= x"0000";
				when 16#1bae# => read_data_o <= x"0000";
				when 16#1baf# => read_data_o <= x"0000";
				when 16#1bb0# => read_data_o <= x"0000";
				when 16#1bb1# => read_data_o <= x"0000";
				when 16#1bb2# => read_data_o <= x"0000";
				when 16#1bb3# => read_data_o <= x"0000";
				when 16#1bb4# => read_data_o <= x"0000";
				when 16#1bb5# => read_data_o <= x"0000";
				when 16#1bb6# => read_data_o <= x"0000";
				when 16#1bb7# => read_data_o <= x"0000";
				when 16#1bb8# => read_data_o <= x"0000";
				when 16#1bb9# => read_data_o <= x"0000";
				when 16#1bba# => read_data_o <= x"0000";
				when 16#1bbb# => read_data_o <= x"0000";
				when 16#1bbc# => read_data_o <= x"0000";
				when 16#1bbd# => read_data_o <= x"0000";
				when 16#1bbe# => read_data_o <= x"0000";
				when 16#1bbf# => read_data_o <= x"0000";
				when 16#1bc0# => read_data_o <= x"0000";
				when 16#1bc1# => read_data_o <= x"0000";
				when 16#1bc2# => read_data_o <= x"0000";
				when 16#1bc3# => read_data_o <= x"0000";
				when 16#1bc4# => read_data_o <= x"0000";
				when 16#1bc5# => read_data_o <= x"0000";
				when 16#1bc6# => read_data_o <= x"0000";
				when 16#1bc7# => read_data_o <= x"0000";
				when 16#1bc8# => read_data_o <= x"0000";
				when 16#1bc9# => read_data_o <= x"0000";
				when 16#1bca# => read_data_o <= x"0000";
				when 16#1bcb# => read_data_o <= x"0000";
				when 16#1bcc# => read_data_o <= x"0000";
				when 16#1bcd# => read_data_o <= x"0000";
				when 16#1bce# => read_data_o <= x"0000";
				when 16#1bcf# => read_data_o <= x"0000";
				when 16#1bd0# => read_data_o <= x"0000";
				when 16#1bd1# => read_data_o <= x"0000";
				when 16#1bd2# => read_data_o <= x"0000";
				when 16#1bd3# => read_data_o <= x"0000";
				when 16#1bd4# => read_data_o <= x"0000";
				when 16#1bd5# => read_data_o <= x"0000";
				when 16#1bd6# => read_data_o <= x"0000";
				when 16#1bd7# => read_data_o <= x"0000";
				when 16#1bd8# => read_data_o <= x"0000";
				when 16#1bd9# => read_data_o <= x"0000";
				when 16#1bda# => read_data_o <= x"0000";
				when 16#1bdb# => read_data_o <= x"0000";
				when 16#1bdc# => read_data_o <= x"0000";
				when 16#1bdd# => read_data_o <= x"0000";
				when 16#1bde# => read_data_o <= x"0000";
				when 16#1bdf# => read_data_o <= x"0000";
				when 16#1be0# => read_data_o <= x"0000";
				when 16#1be1# => read_data_o <= x"0000";
				when 16#1be2# => read_data_o <= x"0000";
				when 16#1be3# => read_data_o <= x"0000";
				when 16#1be4# => read_data_o <= x"0000";
				when 16#1be5# => read_data_o <= x"0000";
				when 16#1be6# => read_data_o <= x"0000";
				when 16#1be7# => read_data_o <= x"0000";
				when 16#1be8# => read_data_o <= x"0000";
				when 16#1be9# => read_data_o <= x"0000";
				when 16#1bea# => read_data_o <= x"0000";
				when 16#1beb# => read_data_o <= x"0000";
				when 16#1bec# => read_data_o <= x"0000";
				when 16#1bed# => read_data_o <= x"0000";
				when 16#1bee# => read_data_o <= x"0000";
				when 16#1bef# => read_data_o <= x"0000";
				when 16#1bf0# => read_data_o <= x"0000";
				when 16#1bf1# => read_data_o <= x"0000";
				when 16#1bf2# => read_data_o <= x"0000";
				when 16#1bf3# => read_data_o <= x"0000";
				when 16#1bf4# => read_data_o <= x"0000";
				when 16#1bf5# => read_data_o <= x"0000";
				when 16#1bf6# => read_data_o <= x"0000";
				when 16#1bf7# => read_data_o <= x"0000";
				when 16#1bf8# => read_data_o <= x"0000";
				when 16#1bf9# => read_data_o <= x"0000";
				when 16#1bfa# => read_data_o <= x"0000";
				when 16#1bfb# => read_data_o <= x"0000";
				when 16#1bfc# => read_data_o <= x"0000";
				when 16#1bfd# => read_data_o <= x"0000";
				when 16#1bfe# => read_data_o <= x"0000";
				when 16#1bff# => read_data_o <= x"0000";
				when 16#1c00# => read_data_o <= x"0000";
				when 16#1c01# => read_data_o <= x"0000";
				when 16#1c02# => read_data_o <= x"0000";
				when 16#1c03# => read_data_o <= x"0000";
				when 16#1c04# => read_data_o <= x"0000";
				when 16#1c05# => read_data_o <= x"0000";
				when 16#1c06# => read_data_o <= x"0000";
				when 16#1c07# => read_data_o <= x"0000";
				when 16#1c08# => read_data_o <= x"0000";
				when 16#1c09# => read_data_o <= x"0000";
				when 16#1c0a# => read_data_o <= x"0000";
				when 16#1c0b# => read_data_o <= x"0000";
				when 16#1c0c# => read_data_o <= x"0000";
				when 16#1c0d# => read_data_o <= x"0000";
				when 16#1c0e# => read_data_o <= x"0000";
				when 16#1c0f# => read_data_o <= x"0000";
				when 16#1c10# => read_data_o <= x"0000";
				when 16#1c11# => read_data_o <= x"0000";
				when 16#1c12# => read_data_o <= x"0000";
				when 16#1c13# => read_data_o <= x"0000";
				when 16#1c14# => read_data_o <= x"0000";
				when 16#1c15# => read_data_o <= x"0000";
				when 16#1c16# => read_data_o <= x"0000";
				when 16#1c17# => read_data_o <= x"0000";
				when 16#1c18# => read_data_o <= x"0000";
				when 16#1c19# => read_data_o <= x"0000";
				when 16#1c1a# => read_data_o <= x"0000";
				when 16#1c1b# => read_data_o <= x"0000";
				when 16#1c1c# => read_data_o <= x"0000";
				when 16#1c1d# => read_data_o <= x"0000";
				when 16#1c1e# => read_data_o <= x"0000";
				when 16#1c1f# => read_data_o <= x"0000";
				when 16#1c20# => read_data_o <= x"0000";
				when 16#1c21# => read_data_o <= x"0000";
				when 16#1c22# => read_data_o <= x"0000";
				when 16#1c23# => read_data_o <= x"0000";
				when 16#1c24# => read_data_o <= x"0000";
				when 16#1c25# => read_data_o <= x"0000";
				when 16#1c26# => read_data_o <= x"0000";
				when 16#1c27# => read_data_o <= x"0000";
				when 16#1c28# => read_data_o <= x"0000";
				when 16#1c29# => read_data_o <= x"0000";
				when 16#1c2a# => read_data_o <= x"0000";
				when 16#1c2b# => read_data_o <= x"0000";
				when 16#1c2c# => read_data_o <= x"0000";
				when 16#1c2d# => read_data_o <= x"0000";
				when 16#1c2e# => read_data_o <= x"0000";
				when 16#1c2f# => read_data_o <= x"0000";
				when 16#1c30# => read_data_o <= x"0000";
				when 16#1c31# => read_data_o <= x"0000";
				when 16#1c32# => read_data_o <= x"0000";
				when 16#1c33# => read_data_o <= x"0000";
				when 16#1c34# => read_data_o <= x"0000";
				when 16#1c35# => read_data_o <= x"0000";
				when 16#1c36# => read_data_o <= x"0000";
				when 16#1c37# => read_data_o <= x"0000";
				when 16#1c38# => read_data_o <= x"0000";
				when 16#1c39# => read_data_o <= x"0000";
				when 16#1c3a# => read_data_o <= x"0000";
				when 16#1c3b# => read_data_o <= x"0000";
				when 16#1c3c# => read_data_o <= x"0000";
				when 16#1c3d# => read_data_o <= x"0000";
				when 16#1c3e# => read_data_o <= x"0000";
				when 16#1c3f# => read_data_o <= x"0000";
				when 16#1c40# => read_data_o <= x"0000";
				when 16#1c41# => read_data_o <= x"0000";
				when 16#1c42# => read_data_o <= x"0000";
				when 16#1c43# => read_data_o <= x"0000";
				when 16#1c44# => read_data_o <= x"0000";
				when 16#1c45# => read_data_o <= x"0000";
				when 16#1c46# => read_data_o <= x"0000";
				when 16#1c47# => read_data_o <= x"0000";
				when 16#1c48# => read_data_o <= x"0000";
				when 16#1c49# => read_data_o <= x"0000";
				when 16#1c4a# => read_data_o <= x"0000";
				when 16#1c4b# => read_data_o <= x"0000";
				when 16#1c4c# => read_data_o <= x"0000";
				when 16#1c4d# => read_data_o <= x"0000";
				when 16#1c4e# => read_data_o <= x"0000";
				when 16#1c4f# => read_data_o <= x"0000";
				when 16#1c50# => read_data_o <= x"0000";
				when 16#1c51# => read_data_o <= x"0000";
				when 16#1c52# => read_data_o <= x"0000";
				when 16#1c53# => read_data_o <= x"0000";
				when 16#1c54# => read_data_o <= x"0000";
				when 16#1c55# => read_data_o <= x"0000";
				when 16#1c56# => read_data_o <= x"0000";
				when 16#1c57# => read_data_o <= x"0000";
				when 16#1c58# => read_data_o <= x"0000";
				when 16#1c59# => read_data_o <= x"0000";
				when 16#1c5a# => read_data_o <= x"0000";
				when 16#1c5b# => read_data_o <= x"0000";
				when 16#1c5c# => read_data_o <= x"0000";
				when 16#1c5d# => read_data_o <= x"0000";
				when 16#1c5e# => read_data_o <= x"0000";
				when 16#1c5f# => read_data_o <= x"0000";
				when 16#1c60# => read_data_o <= x"0000";
				when 16#1c61# => read_data_o <= x"0000";
				when 16#1c62# => read_data_o <= x"0000";
				when 16#1c63# => read_data_o <= x"0000";
				when 16#1c64# => read_data_o <= x"0000";
				when 16#1c65# => read_data_o <= x"0000";
				when 16#1c66# => read_data_o <= x"0000";
				when 16#1c67# => read_data_o <= x"0000";
				when 16#1c68# => read_data_o <= x"0000";
				when 16#1c69# => read_data_o <= x"0000";
				when 16#1c6a# => read_data_o <= x"0000";
				when 16#1c6b# => read_data_o <= x"0000";
				when 16#1c6c# => read_data_o <= x"0000";
				when 16#1c6d# => read_data_o <= x"0000";
				when 16#1c6e# => read_data_o <= x"0000";
				when 16#1c6f# => read_data_o <= x"0000";
				when 16#1c70# => read_data_o <= x"0000";
				when 16#1c71# => read_data_o <= x"0000";
				when 16#1c72# => read_data_o <= x"0000";
				when 16#1c73# => read_data_o <= x"0000";
				when 16#1c74# => read_data_o <= x"0000";
				when 16#1c75# => read_data_o <= x"0000";
				when 16#1c76# => read_data_o <= x"0000";
				when 16#1c77# => read_data_o <= x"0000";
				when 16#1c78# => read_data_o <= x"0000";
				when 16#1c79# => read_data_o <= x"0000";
				when 16#1c7a# => read_data_o <= x"0000";
				when 16#1c7b# => read_data_o <= x"0000";
				when 16#1c7c# => read_data_o <= x"0000";
				when 16#1c7d# => read_data_o <= x"0000";
				when 16#1c7e# => read_data_o <= x"0000";
				when 16#1c7f# => read_data_o <= x"0000";
				when 16#1c80# => read_data_o <= x"0000";
				when 16#1c81# => read_data_o <= x"0000";
				when 16#1c82# => read_data_o <= x"0000";
				when 16#1c83# => read_data_o <= x"0000";
				when 16#1c84# => read_data_o <= x"0000";
				when 16#1c85# => read_data_o <= x"0000";
				when 16#1c86# => read_data_o <= x"0000";
				when 16#1c87# => read_data_o <= x"0000";
				when 16#1c88# => read_data_o <= x"0000";
				when 16#1c89# => read_data_o <= x"0000";
				when 16#1c8a# => read_data_o <= x"0000";
				when 16#1c8b# => read_data_o <= x"0000";
				when 16#1c8c# => read_data_o <= x"0000";
				when 16#1c8d# => read_data_o <= x"0000";
				when 16#1c8e# => read_data_o <= x"0000";
				when 16#1c8f# => read_data_o <= x"0000";
				when 16#1c90# => read_data_o <= x"0000";
				when 16#1c91# => read_data_o <= x"0000";
				when 16#1c92# => read_data_o <= x"0000";
				when 16#1c93# => read_data_o <= x"0000";
				when 16#1c94# => read_data_o <= x"0000";
				when 16#1c95# => read_data_o <= x"0000";
				when 16#1c96# => read_data_o <= x"0000";
				when 16#1c97# => read_data_o <= x"0000";
				when 16#1c98# => read_data_o <= x"0000";
				when 16#1c99# => read_data_o <= x"0000";
				when 16#1c9a# => read_data_o <= x"0000";
				when 16#1c9b# => read_data_o <= x"0000";
				when 16#1c9c# => read_data_o <= x"0000";
				when 16#1c9d# => read_data_o <= x"0000";
				when 16#1c9e# => read_data_o <= x"0000";
				when 16#1c9f# => read_data_o <= x"0000";
				when 16#1ca0# => read_data_o <= x"0000";
				when 16#1ca1# => read_data_o <= x"0000";
				when 16#1ca2# => read_data_o <= x"0000";
				when 16#1ca3# => read_data_o <= x"0000";
				when 16#1ca4# => read_data_o <= x"0000";
				when 16#1ca5# => read_data_o <= x"0000";
				when 16#1ca6# => read_data_o <= x"0000";
				when 16#1ca7# => read_data_o <= x"0000";
				when 16#1ca8# => read_data_o <= x"0000";
				when 16#1ca9# => read_data_o <= x"0000";
				when 16#1caa# => read_data_o <= x"0000";
				when 16#1cab# => read_data_o <= x"0000";
				when 16#1cac# => read_data_o <= x"0000";
				when 16#1cad# => read_data_o <= x"0000";
				when 16#1cae# => read_data_o <= x"0000";
				when 16#1caf# => read_data_o <= x"0000";
				when 16#1cb0# => read_data_o <= x"0000";
				when 16#1cb1# => read_data_o <= x"0000";
				when 16#1cb2# => read_data_o <= x"0000";
				when 16#1cb3# => read_data_o <= x"0000";
				when 16#1cb4# => read_data_o <= x"0000";
				when 16#1cb5# => read_data_o <= x"0000";
				when 16#1cb6# => read_data_o <= x"0000";
				when 16#1cb7# => read_data_o <= x"0000";
				when 16#1cb8# => read_data_o <= x"0000";
				when 16#1cb9# => read_data_o <= x"0000";
				when 16#1cba# => read_data_o <= x"0000";
				when 16#1cbb# => read_data_o <= x"0000";
				when 16#1cbc# => read_data_o <= x"0000";
				when 16#1cbd# => read_data_o <= x"0000";
				when 16#1cbe# => read_data_o <= x"0000";
				when 16#1cbf# => read_data_o <= x"0000";
				when 16#1cc0# => read_data_o <= x"0000";
				when 16#1cc1# => read_data_o <= x"0000";
				when 16#1cc2# => read_data_o <= x"0000";
				when 16#1cc3# => read_data_o <= x"0000";
				when 16#1cc4# => read_data_o <= x"0000";
				when 16#1cc5# => read_data_o <= x"0000";
				when 16#1cc6# => read_data_o <= x"0000";
				when 16#1cc7# => read_data_o <= x"0000";
				when 16#1cc8# => read_data_o <= x"0000";
				when 16#1cc9# => read_data_o <= x"0000";
				when 16#1cca# => read_data_o <= x"0000";
				when 16#1ccb# => read_data_o <= x"0000";
				when 16#1ccc# => read_data_o <= x"0000";
				when 16#1ccd# => read_data_o <= x"0000";
				when 16#1cce# => read_data_o <= x"0000";
				when 16#1ccf# => read_data_o <= x"0000";
				when 16#1cd0# => read_data_o <= x"0000";
				when 16#1cd1# => read_data_o <= x"0000";
				when 16#1cd2# => read_data_o <= x"0000";
				when 16#1cd3# => read_data_o <= x"0000";
				when 16#1cd4# => read_data_o <= x"0000";
				when 16#1cd5# => read_data_o <= x"0000";
				when 16#1cd6# => read_data_o <= x"0000";
				when 16#1cd7# => read_data_o <= x"0000";
				when 16#1cd8# => read_data_o <= x"0000";
				when 16#1cd9# => read_data_o <= x"0000";
				when 16#1cda# => read_data_o <= x"0000";
				when 16#1cdb# => read_data_o <= x"0000";
				when 16#1cdc# => read_data_o <= x"0000";
				when 16#1cdd# => read_data_o <= x"0000";
				when 16#1cde# => read_data_o <= x"0000";
				when 16#1cdf# => read_data_o <= x"0000";
				when 16#1ce0# => read_data_o <= x"0000";
				when 16#1ce1# => read_data_o <= x"0000";
				when 16#1ce2# => read_data_o <= x"0000";
				when 16#1ce3# => read_data_o <= x"0000";
				when 16#1ce4# => read_data_o <= x"0000";
				when 16#1ce5# => read_data_o <= x"0000";
				when 16#1ce6# => read_data_o <= x"0000";
				when 16#1ce7# => read_data_o <= x"0000";
				when 16#1ce8# => read_data_o <= x"0000";
				when 16#1ce9# => read_data_o <= x"0000";
				when 16#1cea# => read_data_o <= x"0000";
				when 16#1ceb# => read_data_o <= x"0000";
				when 16#1cec# => read_data_o <= x"0000";
				when 16#1ced# => read_data_o <= x"0000";
				when 16#1cee# => read_data_o <= x"0000";
				when 16#1cef# => read_data_o <= x"0000";
				when 16#1cf0# => read_data_o <= x"0000";
				when 16#1cf1# => read_data_o <= x"0000";
				when 16#1cf2# => read_data_o <= x"0000";
				when 16#1cf3# => read_data_o <= x"0000";
				when 16#1cf4# => read_data_o <= x"0000";
				when 16#1cf5# => read_data_o <= x"0000";
				when 16#1cf6# => read_data_o <= x"0000";
				when 16#1cf7# => read_data_o <= x"0000";
				when 16#1cf8# => read_data_o <= x"0000";
				when 16#1cf9# => read_data_o <= x"0000";
				when 16#1cfa# => read_data_o <= x"0000";
				when 16#1cfb# => read_data_o <= x"0000";
				when 16#1cfc# => read_data_o <= x"0000";
				when 16#1cfd# => read_data_o <= x"0000";
				when 16#1cfe# => read_data_o <= x"0000";
				when 16#1cff# => read_data_o <= x"0000";
				when 16#1d00# => read_data_o <= x"0000";
				when 16#1d01# => read_data_o <= x"0000";
				when 16#1d02# => read_data_o <= x"0000";
				when 16#1d03# => read_data_o <= x"0000";
				when 16#1d04# => read_data_o <= x"0000";
				when 16#1d05# => read_data_o <= x"0000";
				when 16#1d06# => read_data_o <= x"0000";
				when 16#1d07# => read_data_o <= x"0000";
				when 16#1d08# => read_data_o <= x"0000";
				when 16#1d09# => read_data_o <= x"0000";
				when 16#1d0a# => read_data_o <= x"0000";
				when 16#1d0b# => read_data_o <= x"0000";
				when 16#1d0c# => read_data_o <= x"0000";
				when 16#1d0d# => read_data_o <= x"0000";
				when 16#1d0e# => read_data_o <= x"0000";
				when 16#1d0f# => read_data_o <= x"0000";
				when 16#1d10# => read_data_o <= x"0000";
				when 16#1d11# => read_data_o <= x"0000";
				when 16#1d12# => read_data_o <= x"0000";
				when 16#1d13# => read_data_o <= x"0000";
				when 16#1d14# => read_data_o <= x"0000";
				when 16#1d15# => read_data_o <= x"0000";
				when 16#1d16# => read_data_o <= x"0000";
				when 16#1d17# => read_data_o <= x"0000";
				when 16#1d18# => read_data_o <= x"0000";
				when 16#1d19# => read_data_o <= x"0000";
				when 16#1d1a# => read_data_o <= x"0000";
				when 16#1d1b# => read_data_o <= x"0000";
				when 16#1d1c# => read_data_o <= x"0000";
				when 16#1d1d# => read_data_o <= x"0000";
				when 16#1d1e# => read_data_o <= x"0000";
				when 16#1d1f# => read_data_o <= x"0000";
				when 16#1d20# => read_data_o <= x"0000";
				when 16#1d21# => read_data_o <= x"0000";
				when 16#1d22# => read_data_o <= x"0000";
				when 16#1d23# => read_data_o <= x"0000";
				when 16#1d24# => read_data_o <= x"0000";
				when 16#1d25# => read_data_o <= x"0000";
				when 16#1d26# => read_data_o <= x"0000";
				when 16#1d27# => read_data_o <= x"0000";
				when 16#1d28# => read_data_o <= x"0000";
				when 16#1d29# => read_data_o <= x"0000";
				when 16#1d2a# => read_data_o <= x"0000";
				when 16#1d2b# => read_data_o <= x"0000";
				when 16#1d2c# => read_data_o <= x"0000";
				when 16#1d2d# => read_data_o <= x"0000";
				when 16#1d2e# => read_data_o <= x"0000";
				when 16#1d2f# => read_data_o <= x"0000";
				when 16#1d30# => read_data_o <= x"0000";
				when 16#1d31# => read_data_o <= x"0000";
				when 16#1d32# => read_data_o <= x"0000";
				when 16#1d33# => read_data_o <= x"0000";
				when 16#1d34# => read_data_o <= x"0000";
				when 16#1d35# => read_data_o <= x"0000";
				when 16#1d36# => read_data_o <= x"0000";
				when 16#1d37# => read_data_o <= x"0000";
				when 16#1d38# => read_data_o <= x"0000";
				when 16#1d39# => read_data_o <= x"0000";
				when 16#1d3a# => read_data_o <= x"0000";
				when 16#1d3b# => read_data_o <= x"0000";
				when 16#1d3c# => read_data_o <= x"0000";
				when 16#1d3d# => read_data_o <= x"0000";
				when 16#1d3e# => read_data_o <= x"0000";
				when 16#1d3f# => read_data_o <= x"0000";
				when 16#1d40# => read_data_o <= x"0000";
				when 16#1d41# => read_data_o <= x"0000";
				when 16#1d42# => read_data_o <= x"0000";
				when 16#1d43# => read_data_o <= x"0000";
				when 16#1d44# => read_data_o <= x"0000";
				when 16#1d45# => read_data_o <= x"0000";
				when 16#1d46# => read_data_o <= x"0000";
				when 16#1d47# => read_data_o <= x"0000";
				when 16#1d48# => read_data_o <= x"0000";
				when 16#1d49# => read_data_o <= x"0000";
				when 16#1d4a# => read_data_o <= x"0000";
				when 16#1d4b# => read_data_o <= x"0000";
				when 16#1d4c# => read_data_o <= x"0000";
				when 16#1d4d# => read_data_o <= x"0000";
				when 16#1d4e# => read_data_o <= x"0000";
				when 16#1d4f# => read_data_o <= x"0000";
				when 16#1d50# => read_data_o <= x"0000";
				when 16#1d51# => read_data_o <= x"0000";
				when 16#1d52# => read_data_o <= x"0000";
				when 16#1d53# => read_data_o <= x"0000";
				when 16#1d54# => read_data_o <= x"0000";
				when 16#1d55# => read_data_o <= x"0000";
				when 16#1d56# => read_data_o <= x"0000";
				when 16#1d57# => read_data_o <= x"0000";
				when 16#1d58# => read_data_o <= x"0000";
				when 16#1d59# => read_data_o <= x"0000";
				when 16#1d5a# => read_data_o <= x"0000";
				when 16#1d5b# => read_data_o <= x"0000";
				when 16#1d5c# => read_data_o <= x"0000";
				when 16#1d5d# => read_data_o <= x"0000";
				when 16#1d5e# => read_data_o <= x"0000";
				when 16#1d5f# => read_data_o <= x"0000";
				when 16#1d60# => read_data_o <= x"0000";
				when 16#1d61# => read_data_o <= x"0000";
				when 16#1d62# => read_data_o <= x"0000";
				when 16#1d63# => read_data_o <= x"0000";
				when 16#1d64# => read_data_o <= x"0000";
				when 16#1d65# => read_data_o <= x"0000";
				when 16#1d66# => read_data_o <= x"0000";
				when 16#1d67# => read_data_o <= x"0000";
				when 16#1d68# => read_data_o <= x"0000";
				when 16#1d69# => read_data_o <= x"0000";
				when 16#1d6a# => read_data_o <= x"0000";
				when 16#1d6b# => read_data_o <= x"0000";
				when 16#1d6c# => read_data_o <= x"0000";
				when 16#1d6d# => read_data_o <= x"0000";
				when 16#1d6e# => read_data_o <= x"0000";
				when 16#1d6f# => read_data_o <= x"0000";
				when 16#1d70# => read_data_o <= x"0000";
				when 16#1d71# => read_data_o <= x"0000";
				when 16#1d72# => read_data_o <= x"0000";
				when 16#1d73# => read_data_o <= x"0000";
				when 16#1d74# => read_data_o <= x"0000";
				when 16#1d75# => read_data_o <= x"0000";
				when 16#1d76# => read_data_o <= x"0000";
				when 16#1d77# => read_data_o <= x"0000";
				when 16#1d78# => read_data_o <= x"0000";
				when 16#1d79# => read_data_o <= x"0000";
				when 16#1d7a# => read_data_o <= x"0000";
				when 16#1d7b# => read_data_o <= x"0000";
				when 16#1d7c# => read_data_o <= x"0000";
				when 16#1d7d# => read_data_o <= x"0000";
				when 16#1d7e# => read_data_o <= x"0000";
				when 16#1d7f# => read_data_o <= x"0000";
				when 16#1d80# => read_data_o <= x"0000";
				when 16#1d81# => read_data_o <= x"0000";
				when 16#1d82# => read_data_o <= x"0000";
				when 16#1d83# => read_data_o <= x"0000";
				when 16#1d84# => read_data_o <= x"0000";
				when 16#1d85# => read_data_o <= x"0000";
				when 16#1d86# => read_data_o <= x"0000";
				when 16#1d87# => read_data_o <= x"0000";
				when 16#1d88# => read_data_o <= x"0000";
				when 16#1d89# => read_data_o <= x"0000";
				when 16#1d8a# => read_data_o <= x"0000";
				when 16#1d8b# => read_data_o <= x"0000";
				when 16#1d8c# => read_data_o <= x"0000";
				when 16#1d8d# => read_data_o <= x"0000";
				when 16#1d8e# => read_data_o <= x"0000";
				when 16#1d8f# => read_data_o <= x"0000";
				when 16#1d90# => read_data_o <= x"0000";
				when 16#1d91# => read_data_o <= x"0000";
				when 16#1d92# => read_data_o <= x"0000";
				when 16#1d93# => read_data_o <= x"0000";
				when 16#1d94# => read_data_o <= x"0000";
				when 16#1d95# => read_data_o <= x"0000";
				when 16#1d96# => read_data_o <= x"0000";
				when 16#1d97# => read_data_o <= x"0000";
				when 16#1d98# => read_data_o <= x"0000";
				when 16#1d99# => read_data_o <= x"0000";
				when 16#1d9a# => read_data_o <= x"0000";
				when 16#1d9b# => read_data_o <= x"0000";
				when 16#1d9c# => read_data_o <= x"0000";
				when 16#1d9d# => read_data_o <= x"0000";
				when 16#1d9e# => read_data_o <= x"0000";
				when 16#1d9f# => read_data_o <= x"0000";
				when 16#1da0# => read_data_o <= x"0000";
				when 16#1da1# => read_data_o <= x"0000";
				when 16#1da2# => read_data_o <= x"0000";
				when 16#1da3# => read_data_o <= x"0000";
				when 16#1da4# => read_data_o <= x"0000";
				when 16#1da5# => read_data_o <= x"0000";
				when 16#1da6# => read_data_o <= x"0000";
				when 16#1da7# => read_data_o <= x"0000";
				when 16#1da8# => read_data_o <= x"0000";
				when 16#1da9# => read_data_o <= x"0000";
				when 16#1daa# => read_data_o <= x"0000";
				when 16#1dab# => read_data_o <= x"0000";
				when 16#1dac# => read_data_o <= x"0000";
				when 16#1dad# => read_data_o <= x"0000";
				when 16#1dae# => read_data_o <= x"0000";
				when 16#1daf# => read_data_o <= x"0000";
				when 16#1db0# => read_data_o <= x"0000";
				when 16#1db1# => read_data_o <= x"0000";
				when 16#1db2# => read_data_o <= x"0000";
				when 16#1db3# => read_data_o <= x"0000";
				when 16#1db4# => read_data_o <= x"0000";
				when 16#1db5# => read_data_o <= x"0000";
				when 16#1db6# => read_data_o <= x"0000";
				when 16#1db7# => read_data_o <= x"0000";
				when 16#1db8# => read_data_o <= x"0000";
				when 16#1db9# => read_data_o <= x"0000";
				when 16#1dba# => read_data_o <= x"0000";
				when 16#1dbb# => read_data_o <= x"0000";
				when 16#1dbc# => read_data_o <= x"0000";
				when 16#1dbd# => read_data_o <= x"0000";
				when 16#1dbe# => read_data_o <= x"0000";
				when 16#1dbf# => read_data_o <= x"0000";
				when 16#1dc0# => read_data_o <= x"0000";
				when 16#1dc1# => read_data_o <= x"0000";
				when 16#1dc2# => read_data_o <= x"0000";
				when 16#1dc3# => read_data_o <= x"0000";
				when 16#1dc4# => read_data_o <= x"0000";
				when 16#1dc5# => read_data_o <= x"0000";
				when 16#1dc6# => read_data_o <= x"0000";
				when 16#1dc7# => read_data_o <= x"0000";
				when 16#1dc8# => read_data_o <= x"0000";
				when 16#1dc9# => read_data_o <= x"0000";
				when 16#1dca# => read_data_o <= x"0000";
				when 16#1dcb# => read_data_o <= x"0000";
				when 16#1dcc# => read_data_o <= x"0000";
				when 16#1dcd# => read_data_o <= x"0000";
				when 16#1dce# => read_data_o <= x"0000";
				when 16#1dcf# => read_data_o <= x"0000";
				when 16#1dd0# => read_data_o <= x"0000";
				when 16#1dd1# => read_data_o <= x"0000";
				when 16#1dd2# => read_data_o <= x"0000";
				when 16#1dd3# => read_data_o <= x"0000";
				when 16#1dd4# => read_data_o <= x"0000";
				when 16#1dd5# => read_data_o <= x"0000";
				when 16#1dd6# => read_data_o <= x"0000";
				when 16#1dd7# => read_data_o <= x"0000";
				when 16#1dd8# => read_data_o <= x"0000";
				when 16#1dd9# => read_data_o <= x"0000";
				when 16#1dda# => read_data_o <= x"0000";
				when 16#1ddb# => read_data_o <= x"0000";
				when 16#1ddc# => read_data_o <= x"0000";
				when 16#1ddd# => read_data_o <= x"0000";
				when 16#1dde# => read_data_o <= x"0000";
				when 16#1ddf# => read_data_o <= x"0000";
				when 16#1de0# => read_data_o <= x"0000";
				when 16#1de1# => read_data_o <= x"0000";
				when 16#1de2# => read_data_o <= x"0000";
				when 16#1de3# => read_data_o <= x"0000";
				when 16#1de4# => read_data_o <= x"0000";
				when 16#1de5# => read_data_o <= x"0000";
				when 16#1de6# => read_data_o <= x"0000";
				when 16#1de7# => read_data_o <= x"0000";
				when 16#1de8# => read_data_o <= x"0000";
				when 16#1de9# => read_data_o <= x"0000";
				when 16#1dea# => read_data_o <= x"0000";
				when 16#1deb# => read_data_o <= x"0000";
				when 16#1dec# => read_data_o <= x"0000";
				when 16#1ded# => read_data_o <= x"0000";
				when 16#1dee# => read_data_o <= x"0000";
				when 16#1def# => read_data_o <= x"0000";
				when 16#1df0# => read_data_o <= x"0000";
				when 16#1df1# => read_data_o <= x"0000";
				when 16#1df2# => read_data_o <= x"0000";
				when 16#1df3# => read_data_o <= x"0000";
				when 16#1df4# => read_data_o <= x"0000";
				when 16#1df5# => read_data_o <= x"0000";
				when 16#1df6# => read_data_o <= x"0000";
				when 16#1df7# => read_data_o <= x"0000";
				when 16#1df8# => read_data_o <= x"0000";
				when 16#1df9# => read_data_o <= x"0000";
				when 16#1dfa# => read_data_o <= x"0000";
				when 16#1dfb# => read_data_o <= x"0000";
				when 16#1dfc# => read_data_o <= x"0000";
				when 16#1dfd# => read_data_o <= x"0000";
				when 16#1dfe# => read_data_o <= x"0000";
				when 16#1dff# => read_data_o <= x"0000";
				when 16#1e00# => read_data_o <= x"0000";
				when 16#1e01# => read_data_o <= x"0000";
				when 16#1e02# => read_data_o <= x"0000";
				when 16#1e03# => read_data_o <= x"0000";
				when 16#1e04# => read_data_o <= x"0000";
				when 16#1e05# => read_data_o <= x"0000";
				when 16#1e06# => read_data_o <= x"0000";
				when 16#1e07# => read_data_o <= x"0000";
				when 16#1e08# => read_data_o <= x"0000";
				when 16#1e09# => read_data_o <= x"0000";
				when 16#1e0a# => read_data_o <= x"0000";
				when 16#1e0b# => read_data_o <= x"0000";
				when 16#1e0c# => read_data_o <= x"0000";
				when 16#1e0d# => read_data_o <= x"0000";
				when 16#1e0e# => read_data_o <= x"0000";
				when 16#1e0f# => read_data_o <= x"0000";
				when 16#1e10# => read_data_o <= x"0000";
				when 16#1e11# => read_data_o <= x"0000";
				when 16#1e12# => read_data_o <= x"0000";
				when 16#1e13# => read_data_o <= x"0000";
				when 16#1e14# => read_data_o <= x"0000";
				when 16#1e15# => read_data_o <= x"0000";
				when 16#1e16# => read_data_o <= x"0000";
				when 16#1e17# => read_data_o <= x"0000";
				when 16#1e18# => read_data_o <= x"0000";
				when 16#1e19# => read_data_o <= x"0000";
				when 16#1e1a# => read_data_o <= x"0000";
				when 16#1e1b# => read_data_o <= x"0000";
				when 16#1e1c# => read_data_o <= x"0000";
				when 16#1e1d# => read_data_o <= x"0000";
				when 16#1e1e# => read_data_o <= x"0000";
				when 16#1e1f# => read_data_o <= x"0000";
				when 16#1e20# => read_data_o <= x"0000";
				when 16#1e21# => read_data_o <= x"0000";
				when 16#1e22# => read_data_o <= x"0000";
				when 16#1e23# => read_data_o <= x"0000";
				when 16#1e24# => read_data_o <= x"0000";
				when 16#1e25# => read_data_o <= x"0000";
				when 16#1e26# => read_data_o <= x"0000";
				when 16#1e27# => read_data_o <= x"0000";
				when 16#1e28# => read_data_o <= x"0000";
				when 16#1e29# => read_data_o <= x"0000";
				when 16#1e2a# => read_data_o <= x"0000";
				when 16#1e2b# => read_data_o <= x"0000";
				when 16#1e2c# => read_data_o <= x"0000";
				when 16#1e2d# => read_data_o <= x"0000";
				when 16#1e2e# => read_data_o <= x"0000";
				when 16#1e2f# => read_data_o <= x"0000";
				when 16#1e30# => read_data_o <= x"0000";
				when 16#1e31# => read_data_o <= x"0000";
				when 16#1e32# => read_data_o <= x"0000";
				when 16#1e33# => read_data_o <= x"0000";
				when 16#1e34# => read_data_o <= x"0000";
				when 16#1e35# => read_data_o <= x"0000";
				when 16#1e36# => read_data_o <= x"0000";
				when 16#1e37# => read_data_o <= x"0000";
				when 16#1e38# => read_data_o <= x"0000";
				when 16#1e39# => read_data_o <= x"0000";
				when 16#1e3a# => read_data_o <= x"0000";
				when 16#1e3b# => read_data_o <= x"0000";
				when 16#1e3c# => read_data_o <= x"0000";
				when 16#1e3d# => read_data_o <= x"0000";
				when 16#1e3e# => read_data_o <= x"0000";
				when 16#1e3f# => read_data_o <= x"0000";
				when 16#1e40# => read_data_o <= x"0000";
				when 16#1e41# => read_data_o <= x"0000";
				when 16#1e42# => read_data_o <= x"0000";
				when 16#1e43# => read_data_o <= x"0000";
				when 16#1e44# => read_data_o <= x"0000";
				when 16#1e45# => read_data_o <= x"0000";
				when 16#1e46# => read_data_o <= x"0000";
				when 16#1e47# => read_data_o <= x"0000";
				when 16#1e48# => read_data_o <= x"0000";
				when 16#1e49# => read_data_o <= x"0000";
				when 16#1e4a# => read_data_o <= x"0000";
				when 16#1e4b# => read_data_o <= x"0000";
				when 16#1e4c# => read_data_o <= x"0000";
				when 16#1e4d# => read_data_o <= x"0000";
				when 16#1e4e# => read_data_o <= x"0000";
				when 16#1e4f# => read_data_o <= x"0000";
				when 16#1e50# => read_data_o <= x"0000";
				when 16#1e51# => read_data_o <= x"0000";
				when 16#1e52# => read_data_o <= x"0000";
				when 16#1e53# => read_data_o <= x"0000";
				when 16#1e54# => read_data_o <= x"0000";
				when 16#1e55# => read_data_o <= x"0000";
				when 16#1e56# => read_data_o <= x"0000";
				when 16#1e57# => read_data_o <= x"0000";
				when 16#1e58# => read_data_o <= x"0000";
				when 16#1e59# => read_data_o <= x"0000";
				when 16#1e5a# => read_data_o <= x"0000";
				when 16#1e5b# => read_data_o <= x"0000";
				when 16#1e5c# => read_data_o <= x"0000";
				when 16#1e5d# => read_data_o <= x"0000";
				when 16#1e5e# => read_data_o <= x"0000";
				when 16#1e5f# => read_data_o <= x"0000";
				when 16#1e60# => read_data_o <= x"0000";
				when 16#1e61# => read_data_o <= x"0000";
				when 16#1e62# => read_data_o <= x"0000";
				when 16#1e63# => read_data_o <= x"0000";
				when 16#1e64# => read_data_o <= x"0000";
				when 16#1e65# => read_data_o <= x"0000";
				when 16#1e66# => read_data_o <= x"0000";
				when 16#1e67# => read_data_o <= x"0000";
				when 16#1e68# => read_data_o <= x"0000";
				when 16#1e69# => read_data_o <= x"0000";
				when 16#1e6a# => read_data_o <= x"0000";
				when 16#1e6b# => read_data_o <= x"0000";
				when 16#1e6c# => read_data_o <= x"0000";
				when 16#1e6d# => read_data_o <= x"0000";
				when 16#1e6e# => read_data_o <= x"0000";
				when 16#1e6f# => read_data_o <= x"0000";
				when 16#1e70# => read_data_o <= x"0000";
				when 16#1e71# => read_data_o <= x"0000";
				when 16#1e72# => read_data_o <= x"0000";
				when 16#1e73# => read_data_o <= x"0000";
				when 16#1e74# => read_data_o <= x"0000";
				when 16#1e75# => read_data_o <= x"0000";
				when 16#1e76# => read_data_o <= x"0000";
				when 16#1e77# => read_data_o <= x"0000";
				when 16#1e78# => read_data_o <= x"0000";
				when 16#1e79# => read_data_o <= x"0000";
				when 16#1e7a# => read_data_o <= x"0000";
				when 16#1e7b# => read_data_o <= x"0000";
				when 16#1e7c# => read_data_o <= x"0000";
				when 16#1e7d# => read_data_o <= x"0000";
				when 16#1e7e# => read_data_o <= x"0000";
				when 16#1e7f# => read_data_o <= x"0000";
				when 16#1e80# => read_data_o <= x"0000";
				when 16#1e81# => read_data_o <= x"0000";
				when 16#1e82# => read_data_o <= x"0000";
				when 16#1e83# => read_data_o <= x"0000";
				when 16#1e84# => read_data_o <= x"0000";
				when 16#1e85# => read_data_o <= x"0000";
				when 16#1e86# => read_data_o <= x"0000";
				when 16#1e87# => read_data_o <= x"0000";
				when 16#1e88# => read_data_o <= x"0000";
				when 16#1e89# => read_data_o <= x"0000";
				when 16#1e8a# => read_data_o <= x"0000";
				when 16#1e8b# => read_data_o <= x"0000";
				when 16#1e8c# => read_data_o <= x"0000";
				when 16#1e8d# => read_data_o <= x"0000";
				when 16#1e8e# => read_data_o <= x"0000";
				when 16#1e8f# => read_data_o <= x"0000";
				when 16#1e90# => read_data_o <= x"0000";
				when 16#1e91# => read_data_o <= x"0000";
				when 16#1e92# => read_data_o <= x"0000";
				when 16#1e93# => read_data_o <= x"0000";
				when 16#1e94# => read_data_o <= x"0000";
				when 16#1e95# => read_data_o <= x"0000";
				when 16#1e96# => read_data_o <= x"0000";
				when 16#1e97# => read_data_o <= x"0000";
				when 16#1e98# => read_data_o <= x"0000";
				when 16#1e99# => read_data_o <= x"0000";
				when 16#1e9a# => read_data_o <= x"0000";
				when 16#1e9b# => read_data_o <= x"0000";
				when 16#1e9c# => read_data_o <= x"0000";
				when 16#1e9d# => read_data_o <= x"0000";
				when 16#1e9e# => read_data_o <= x"0000";
				when 16#1e9f# => read_data_o <= x"0000";
				when 16#1ea0# => read_data_o <= x"0000";
				when 16#1ea1# => read_data_o <= x"0000";
				when 16#1ea2# => read_data_o <= x"0000";
				when 16#1ea3# => read_data_o <= x"0000";
				when 16#1ea4# => read_data_o <= x"0000";
				when 16#1ea5# => read_data_o <= x"0000";
				when 16#1ea6# => read_data_o <= x"0000";
				when 16#1ea7# => read_data_o <= x"0000";
				when 16#1ea8# => read_data_o <= x"0000";
				when 16#1ea9# => read_data_o <= x"0000";
				when 16#1eaa# => read_data_o <= x"0000";
				when 16#1eab# => read_data_o <= x"0000";
				when 16#1eac# => read_data_o <= x"0000";
				when 16#1ead# => read_data_o <= x"0000";
				when 16#1eae# => read_data_o <= x"0000";
				when 16#1eaf# => read_data_o <= x"0000";
				when 16#1eb0# => read_data_o <= x"0000";
				when 16#1eb1# => read_data_o <= x"0000";
				when 16#1eb2# => read_data_o <= x"0000";
				when 16#1eb3# => read_data_o <= x"0000";
				when 16#1eb4# => read_data_o <= x"0000";
				when 16#1eb5# => read_data_o <= x"0000";
				when 16#1eb6# => read_data_o <= x"0000";
				when 16#1eb7# => read_data_o <= x"0000";
				when 16#1eb8# => read_data_o <= x"0000";
				when 16#1eb9# => read_data_o <= x"0000";
				when 16#1eba# => read_data_o <= x"0000";
				when 16#1ebb# => read_data_o <= x"0000";
				when 16#1ebc# => read_data_o <= x"0000";
				when 16#1ebd# => read_data_o <= x"0000";
				when 16#1ebe# => read_data_o <= x"0000";
				when 16#1ebf# => read_data_o <= x"0000";
				when 16#1ec0# => read_data_o <= x"0000";
				when 16#1ec1# => read_data_o <= x"0000";
				when 16#1ec2# => read_data_o <= x"0000";
				when 16#1ec3# => read_data_o <= x"0000";
				when 16#1ec4# => read_data_o <= x"0000";
				when 16#1ec5# => read_data_o <= x"0000";
				when 16#1ec6# => read_data_o <= x"0000";
				when 16#1ec7# => read_data_o <= x"0000";
				when 16#1ec8# => read_data_o <= x"0000";
				when 16#1ec9# => read_data_o <= x"0000";
				when 16#1eca# => read_data_o <= x"0000";
				when 16#1ecb# => read_data_o <= x"0000";
				when 16#1ecc# => read_data_o <= x"0000";
				when 16#1ecd# => read_data_o <= x"0000";
				when 16#1ece# => read_data_o <= x"0000";
				when 16#1ecf# => read_data_o <= x"0000";
				when 16#1ed0# => read_data_o <= x"0000";
				when 16#1ed1# => read_data_o <= x"0000";
				when 16#1ed2# => read_data_o <= x"0000";
				when 16#1ed3# => read_data_o <= x"0000";
				when 16#1ed4# => read_data_o <= x"0000";
				when 16#1ed5# => read_data_o <= x"0000";
				when 16#1ed6# => read_data_o <= x"0000";
				when 16#1ed7# => read_data_o <= x"0000";
				when 16#1ed8# => read_data_o <= x"0000";
				when 16#1ed9# => read_data_o <= x"0000";
				when 16#1eda# => read_data_o <= x"0000";
				when 16#1edb# => read_data_o <= x"0000";
				when 16#1edc# => read_data_o <= x"0000";
				when 16#1edd# => read_data_o <= x"0000";
				when 16#1ede# => read_data_o <= x"0000";
				when 16#1edf# => read_data_o <= x"0000";
				when 16#1ee0# => read_data_o <= x"0000";
				when 16#1ee1# => read_data_o <= x"0000";
				when 16#1ee2# => read_data_o <= x"0000";
				when 16#1ee3# => read_data_o <= x"0000";
				when 16#1ee4# => read_data_o <= x"0000";
				when 16#1ee5# => read_data_o <= x"0000";
				when 16#1ee6# => read_data_o <= x"0000";
				when 16#1ee7# => read_data_o <= x"0000";
				when 16#1ee8# => read_data_o <= x"0000";
				when 16#1ee9# => read_data_o <= x"0000";
				when 16#1eea# => read_data_o <= x"0000";
				when 16#1eeb# => read_data_o <= x"0000";
				when 16#1eec# => read_data_o <= x"0000";
				when 16#1eed# => read_data_o <= x"0000";
				when 16#1eee# => read_data_o <= x"0000";
				when 16#1eef# => read_data_o <= x"0000";
				when 16#1ef0# => read_data_o <= x"0000";
				when 16#1ef1# => read_data_o <= x"0000";
				when 16#1ef2# => read_data_o <= x"0000";
				when 16#1ef3# => read_data_o <= x"0000";
				when 16#1ef4# => read_data_o <= x"0000";
				when 16#1ef5# => read_data_o <= x"0000";
				when 16#1ef6# => read_data_o <= x"0000";
				when 16#1ef7# => read_data_o <= x"0000";
				when 16#1ef8# => read_data_o <= x"0000";
				when 16#1ef9# => read_data_o <= x"0000";
				when 16#1efa# => read_data_o <= x"0000";
				when 16#1efb# => read_data_o <= x"0000";
				when 16#1efc# => read_data_o <= x"0000";
				when 16#1efd# => read_data_o <= x"0000";
				when 16#1efe# => read_data_o <= x"0000";
				when 16#1eff# => read_data_o <= x"0000";
				when 16#1f00# => read_data_o <= x"0000";
				when 16#1f01# => read_data_o <= x"0000";
				when 16#1f02# => read_data_o <= x"0000";
				when 16#1f03# => read_data_o <= x"0000";
				when 16#1f04# => read_data_o <= x"0000";
				when 16#1f05# => read_data_o <= x"0000";
				when 16#1f06# => read_data_o <= x"0000";
				when 16#1f07# => read_data_o <= x"0000";
				when 16#1f08# => read_data_o <= x"0000";
				when 16#1f09# => read_data_o <= x"0000";
				when 16#1f0a# => read_data_o <= x"0000";
				when 16#1f0b# => read_data_o <= x"0000";
				when 16#1f0c# => read_data_o <= x"0000";
				when 16#1f0d# => read_data_o <= x"0000";
				when 16#1f0e# => read_data_o <= x"0000";
				when 16#1f0f# => read_data_o <= x"0000";
				when 16#1f10# => read_data_o <= x"0000";
				when 16#1f11# => read_data_o <= x"0000";
				when 16#1f12# => read_data_o <= x"0000";
				when 16#1f13# => read_data_o <= x"0000";
				when 16#1f14# => read_data_o <= x"0000";
				when 16#1f15# => read_data_o <= x"0000";
				when 16#1f16# => read_data_o <= x"0000";
				when 16#1f17# => read_data_o <= x"0000";
				when 16#1f18# => read_data_o <= x"0000";
				when 16#1f19# => read_data_o <= x"0000";
				when 16#1f1a# => read_data_o <= x"0000";
				when 16#1f1b# => read_data_o <= x"0000";
				when 16#1f1c# => read_data_o <= x"0000";
				when 16#1f1d# => read_data_o <= x"0000";
				when 16#1f1e# => read_data_o <= x"0000";
				when 16#1f1f# => read_data_o <= x"0000";
				when 16#1f20# => read_data_o <= x"0000";
				when 16#1f21# => read_data_o <= x"0000";
				when 16#1f22# => read_data_o <= x"0000";
				when 16#1f23# => read_data_o <= x"0000";
				when 16#1f24# => read_data_o <= x"0000";
				when 16#1f25# => read_data_o <= x"0000";
				when 16#1f26# => read_data_o <= x"0000";
				when 16#1f27# => read_data_o <= x"0000";
				when 16#1f28# => read_data_o <= x"0000";
				when 16#1f29# => read_data_o <= x"0000";
				when 16#1f2a# => read_data_o <= x"0000";
				when 16#1f2b# => read_data_o <= x"0000";
				when 16#1f2c# => read_data_o <= x"0000";
				when 16#1f2d# => read_data_o <= x"0000";
				when 16#1f2e# => read_data_o <= x"0000";
				when 16#1f2f# => read_data_o <= x"0000";
				when 16#1f30# => read_data_o <= x"0000";
				when 16#1f31# => read_data_o <= x"0000";
				when 16#1f32# => read_data_o <= x"0000";
				when 16#1f33# => read_data_o <= x"0000";
				when 16#1f34# => read_data_o <= x"0000";
				when 16#1f35# => read_data_o <= x"0000";
				when 16#1f36# => read_data_o <= x"0000";
				when 16#1f37# => read_data_o <= x"0000";
				when 16#1f38# => read_data_o <= x"0000";
				when 16#1f39# => read_data_o <= x"0000";
				when 16#1f3a# => read_data_o <= x"0000";
				when 16#1f3b# => read_data_o <= x"0000";
				when 16#1f3c# => read_data_o <= x"0000";
				when 16#1f3d# => read_data_o <= x"0000";
				when 16#1f3e# => read_data_o <= x"0000";
				when 16#1f3f# => read_data_o <= x"0000";
				when 16#1f40# => read_data_o <= x"0000";
				when 16#1f41# => read_data_o <= x"0000";
				when 16#1f42# => read_data_o <= x"0000";
				when 16#1f43# => read_data_o <= x"0000";
				when 16#1f44# => read_data_o <= x"0000";
				when 16#1f45# => read_data_o <= x"0000";
				when 16#1f46# => read_data_o <= x"0000";
				when 16#1f47# => read_data_o <= x"0000";
				when 16#1f48# => read_data_o <= x"0000";
				when 16#1f49# => read_data_o <= x"0000";
				when 16#1f4a# => read_data_o <= x"0000";
				when 16#1f4b# => read_data_o <= x"0000";
				when 16#1f4c# => read_data_o <= x"0000";
				when 16#1f4d# => read_data_o <= x"0000";
				when 16#1f4e# => read_data_o <= x"0000";
				when 16#1f4f# => read_data_o <= x"0000";
				when 16#1f50# => read_data_o <= x"0000";
				when 16#1f51# => read_data_o <= x"0000";
				when 16#1f52# => read_data_o <= x"0000";
				when 16#1f53# => read_data_o <= x"0000";
				when 16#1f54# => read_data_o <= x"0000";
				when 16#1f55# => read_data_o <= x"0000";
				when 16#1f56# => read_data_o <= x"0000";
				when 16#1f57# => read_data_o <= x"0000";
				when 16#1f58# => read_data_o <= x"0000";
				when 16#1f59# => read_data_o <= x"0000";
				when 16#1f5a# => read_data_o <= x"0000";
				when 16#1f5b# => read_data_o <= x"0000";
				when 16#1f5c# => read_data_o <= x"0000";
				when 16#1f5d# => read_data_o <= x"0000";
				when 16#1f5e# => read_data_o <= x"0000";
				when 16#1f5f# => read_data_o <= x"0000";
				when 16#1f60# => read_data_o <= x"0000";
				when 16#1f61# => read_data_o <= x"0000";
				when 16#1f62# => read_data_o <= x"0000";
				when 16#1f63# => read_data_o <= x"0000";
				when 16#1f64# => read_data_o <= x"0000";
				when 16#1f65# => read_data_o <= x"0000";
				when 16#1f66# => read_data_o <= x"0000";
				when 16#1f67# => read_data_o <= x"0000";
				when 16#1f68# => read_data_o <= x"0000";
				when 16#1f69# => read_data_o <= x"0000";
				when 16#1f6a# => read_data_o <= x"0000";
				when 16#1f6b# => read_data_o <= x"0000";
				when 16#1f6c# => read_data_o <= x"0000";
				when 16#1f6d# => read_data_o <= x"0000";
				when 16#1f6e# => read_data_o <= x"0000";
				when 16#1f6f# => read_data_o <= x"0000";
				when 16#1f70# => read_data_o <= x"0000";
				when 16#1f71# => read_data_o <= x"0000";
				when 16#1f72# => read_data_o <= x"0000";
				when 16#1f73# => read_data_o <= x"0000";
				when 16#1f74# => read_data_o <= x"0000";
				when 16#1f75# => read_data_o <= x"0000";
				when 16#1f76# => read_data_o <= x"0000";
				when 16#1f77# => read_data_o <= x"0000";
				when 16#1f78# => read_data_o <= x"0000";
				when 16#1f79# => read_data_o <= x"0000";
				when 16#1f7a# => read_data_o <= x"0000";
				when 16#1f7b# => read_data_o <= x"0000";
				when 16#1f7c# => read_data_o <= x"0000";
				when 16#1f7d# => read_data_o <= x"0000";
				when 16#1f7e# => read_data_o <= x"0000";
				when 16#1f7f# => read_data_o <= x"0000";
				when 16#1f80# => read_data_o <= x"0000";
				when 16#1f81# => read_data_o <= x"0000";
				when 16#1f82# => read_data_o <= x"0000";
				when 16#1f83# => read_data_o <= x"0000";
				when 16#1f84# => read_data_o <= x"0000";
				when 16#1f85# => read_data_o <= x"0000";
				when 16#1f86# => read_data_o <= x"0000";
				when 16#1f87# => read_data_o <= x"0000";
				when 16#1f88# => read_data_o <= x"0000";
				when 16#1f89# => read_data_o <= x"0000";
				when 16#1f8a# => read_data_o <= x"0000";
				when 16#1f8b# => read_data_o <= x"0000";
				when 16#1f8c# => read_data_o <= x"0000";
				when 16#1f8d# => read_data_o <= x"0000";
				when 16#1f8e# => read_data_o <= x"0000";
				when 16#1f8f# => read_data_o <= x"0000";
				when 16#1f90# => read_data_o <= x"0000";
				when 16#1f91# => read_data_o <= x"0000";
				when 16#1f92# => read_data_o <= x"0000";
				when 16#1f93# => read_data_o <= x"0000";
				when 16#1f94# => read_data_o <= x"0000";
				when 16#1f95# => read_data_o <= x"0000";
				when 16#1f96# => read_data_o <= x"0000";
				when 16#1f97# => read_data_o <= x"0000";
				when 16#1f98# => read_data_o <= x"0000";
				when 16#1f99# => read_data_o <= x"0000";
				when 16#1f9a# => read_data_o <= x"0000";
				when 16#1f9b# => read_data_o <= x"0000";
				when 16#1f9c# => read_data_o <= x"0000";
				when 16#1f9d# => read_data_o <= x"0000";
				when 16#1f9e# => read_data_o <= x"0000";
				when 16#1f9f# => read_data_o <= x"0000";
				when 16#1fa0# => read_data_o <= x"0000";
				when 16#1fa1# => read_data_o <= x"0000";
				when 16#1fa2# => read_data_o <= x"0000";
				when 16#1fa3# => read_data_o <= x"0000";
				when 16#1fa4# => read_data_o <= x"0000";
				when 16#1fa5# => read_data_o <= x"0000";
				when 16#1fa6# => read_data_o <= x"0000";
				when 16#1fa7# => read_data_o <= x"0000";
				when 16#1fa8# => read_data_o <= x"0000";
				when 16#1fa9# => read_data_o <= x"0000";
				when 16#1faa# => read_data_o <= x"0000";
				when 16#1fab# => read_data_o <= x"0000";
				when 16#1fac# => read_data_o <= x"0000";
				when 16#1fad# => read_data_o <= x"0000";
				when 16#1fae# => read_data_o <= x"0000";
				when 16#1faf# => read_data_o <= x"0000";
				when 16#1fb0# => read_data_o <= x"0000";
				when 16#1fb1# => read_data_o <= x"0000";
				when 16#1fb2# => read_data_o <= x"0000";
				when 16#1fb3# => read_data_o <= x"0000";
				when 16#1fb4# => read_data_o <= x"0000";
				when 16#1fb5# => read_data_o <= x"0000";
				when 16#1fb6# => read_data_o <= x"0000";
				when 16#1fb7# => read_data_o <= x"0000";
				when 16#1fb8# => read_data_o <= x"0000";
				when 16#1fb9# => read_data_o <= x"0000";
				when 16#1fba# => read_data_o <= x"0000";
				when 16#1fbb# => read_data_o <= x"0000";
				when 16#1fbc# => read_data_o <= x"0000";
				when 16#1fbd# => read_data_o <= x"0000";
				when 16#1fbe# => read_data_o <= x"0000";
				when 16#1fbf# => read_data_o <= x"0000";
				when 16#1fc0# => read_data_o <= x"0000";
				when 16#1fc1# => read_data_o <= x"0000";
				when 16#1fc2# => read_data_o <= x"0000";
				when 16#1fc3# => read_data_o <= x"0000";
				when 16#1fc4# => read_data_o <= x"0000";
				when 16#1fc5# => read_data_o <= x"0000";
				when 16#1fc6# => read_data_o <= x"0000";
				when 16#1fc7# => read_data_o <= x"0000";
				when 16#1fc8# => read_data_o <= x"0000";
				when 16#1fc9# => read_data_o <= x"0000";
				when 16#1fca# => read_data_o <= x"0000";
				when 16#1fcb# => read_data_o <= x"0000";
				when 16#1fcc# => read_data_o <= x"0000";
				when 16#1fcd# => read_data_o <= x"0000";
				when 16#1fce# => read_data_o <= x"0000";
				when 16#1fcf# => read_data_o <= x"0000";
				when 16#1fd0# => read_data_o <= x"0000";
				when 16#1fd1# => read_data_o <= x"0000";
				when 16#1fd2# => read_data_o <= x"0000";
				when 16#1fd3# => read_data_o <= x"0000";
				when 16#1fd4# => read_data_o <= x"0000";
				when 16#1fd5# => read_data_o <= x"0000";
				when 16#1fd6# => read_data_o <= x"0000";
				when 16#1fd7# => read_data_o <= x"0000";
				when 16#1fd8# => read_data_o <= x"0000";
				when 16#1fd9# => read_data_o <= x"0000";
				when 16#1fda# => read_data_o <= x"0000";
				when 16#1fdb# => read_data_o <= x"0000";
				when 16#1fdc# => read_data_o <= x"0000";
				when 16#1fdd# => read_data_o <= x"0000";
				when 16#1fde# => read_data_o <= x"0000";
				when 16#1fdf# => read_data_o <= x"0000";
				when 16#1fe0# => read_data_o <= x"0000";
				when 16#1fe1# => read_data_o <= x"0000";
				when 16#1fe2# => read_data_o <= x"0000";
				when 16#1fe3# => read_data_o <= x"0000";
				when 16#1fe4# => read_data_o <= x"0000";
				when 16#1fe5# => read_data_o <= x"0000";
				when 16#1fe6# => read_data_o <= x"0000";
				when 16#1fe7# => read_data_o <= x"0000";
				when 16#1fe8# => read_data_o <= x"0000";
				when 16#1fe9# => read_data_o <= x"0000";
				when 16#1fea# => read_data_o <= x"0000";
				when 16#1feb# => read_data_o <= x"0000";
				when 16#1fec# => read_data_o <= x"0000";
				when 16#1fed# => read_data_o <= x"0000";
				when 16#1fee# => read_data_o <= x"0000";
				when 16#1fef# => read_data_o <= x"0000";
				when 16#1ff0# => read_data_o <= x"0000";
				when 16#1ff1# => read_data_o <= x"0000";
				when 16#1ff2# => read_data_o <= x"0000";
				when 16#1ff3# => read_data_o <= x"0000";
				when 16#1ff4# => read_data_o <= x"0000";
				when 16#1ff5# => read_data_o <= x"0000";
				when 16#1ff6# => read_data_o <= x"0000";
				when 16#1ff7# => read_data_o <= x"0000";
				when 16#1ff8# => read_data_o <= x"0000";
				when 16#1ff9# => read_data_o <= x"0000";
				when 16#1ffa# => read_data_o <= x"0000";
				when 16#1ffb# => read_data_o <= x"0000";
				when 16#1ffc# => read_data_o <= x"0000";
				when 16#1ffd# => read_data_o <= x"0000";
				when 16#1ffe# => read_data_o <= x"0000";
				when 16#1fff# => read_data_o <= x"0000";
				when others => read_data_o <= x"a000";
			end case;
		end if;
	end process;

end rtl;
