library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library unisim;
use unisim.Vcomponents.all;
library unimacro;
use unimacro.Vcomponents.all;
entity fontrom is port(
	clk_i  : in std_logic;
	addr_i : in integer;
	data_o : out std_logic_vector(0 downto 0));
end fontrom;

architecture rtl of fontrom is

signal rom_addr_s: std_logic_vector(15 downto 0);
signal rom_data_s: std_logic_vector(31 downto 0);
signal data0_s: std_logic_vector(0 downto 0);
signal data1_s: std_logic_vector(0 downto 0);
signal data2_s: std_logic_vector(0 downto 0);
begin

	rom0: RAMB16_S1
		generic map(
			INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0008006001800600180060000000000000000000000000000000000000000000",
INIT_16 => X"00000000000000000000000000000000000CC066019800000000180060000002",
INIT_17 => X"36007E006C199836C07E0060000019806607FE1FF819806607FE1FF819806600",
INIT_18 => X"000000000000E186CC1B603B001800DC06D83361870000000006007E036C1998",
INIT_19 => X"00000000000001C00C003800E000001C06CC0E182CC1160070036018C0760070",
INIT_1A => X"18003800001C0018003000600180060018006003001801C00000000000000000",
INIT_1B => X"199876E03C00F01DB86660180060000003801800C00600180060018006000C00",
INIT_1C => X"000000000000000018006001803FC0FF00600180060000000000000000180060",
INIT_1D => X"000000FFF3FFC00000000000000000000007003000E000000000000000000000",
INIT_1E => X"6003000800000000003800E00000000000000000000000000000000000000000",
INIT_1F => X"01980C3030C0C3030C0C3030C06600F0000C006003001800C006003001800C00",
INIT_20 => X"006060C301F800000000FF006001800600180060019007801C0060000000003C",
INIT_21 => X"7E030C18186000C001F00C006060C301F800000001FF80060070070070030018",
INIT_22 => X"07F800600183FE000000006001801FF8186063019806C01E0070018000000000",
INIT_23 => X"007E030C18186060C381F6001800C0C601F0000000007E030C18186001800300",
INIT_24 => X"F80C306060C301F80000000006001800C006003001800C0060018007FE000000",
INIT_25 => X"00003E018C0C006001BE070C18186060C301F8000000007E030C18186060C301",
INIT_26 => X"00E000000000000000000000003800E0000000003800E0000000000000000000",
INIT_27 => X"00080030006000C0018006003001800C00200000000007003000E00000000038",
INIT_28 => X"6000C001800300040000000000000003FC0FF000000003FC0FF0000000000000",
INIT_29 => X"000000003800E000000E0030038018006060C301F8000001000C006003001800",
INIT_2A => X"C0C3030C066019803C00F00001FE07FC00387E61F987E61F9830E0FF01F80000",
INIT_2B => X"F0000000007F830618186060C181FE0C186060C181FE0000000181860618183F",
INIT_2C => X"6061818606181830606180FE000000007C031818300060018006001860C0C601",
INIT_2D => X"87FE00000001FF8006001800600181FE001800600187FE000000003F81860C18",
INIT_2E => X"306061F18006001860C0C601F000000000018006001800607F80060018006001",
INIT_2F => X"1801F800000001818606181860618187FE1818606181860600000001BC071818",
INIT_30 => X"0C006001800600180060018007F0000000007E00600180060018006001800600",
INIT_31 => X"60018006000000018186060C18186031807E03181860C18606000000003F0186",
INIT_32 => X"06181860619986F61E7870E181840200000001FF800600180060018006001800",
INIT_33 => X"30C06600F0000000018186061C187861B1866618D861E1838606000000018186",
INIT_34 => X"8006001800607F830618186060C181FE000000003C01980C3060618186061818",
INIT_35 => X"186060C181FE0C0038003C01D80DB06061818606181830C06600F00000000001",
INIT_36 => X"7E030C18186000C001F800300060C301F8000000018186060C1818607F830618",
INIT_37 => X"181860618186060000000018006001800600180060018006001807FE00000000",
INIT_38 => X"003C00F006601980C3030C0C306061818606000000003C01980C306061818606",
INIT_39 => X"6003C01980C30606000000006601980FF036C0DB066619986061818606000000",
INIT_3A => X"0000180060018006001800F0066030C1818606000000018186060C3019803C00",
INIT_3B => X"0018006001800601F800000001FF800C006003001800C0060030018007FE0000",
INIT_3C => X"006000C00180030006000C00180030006000C00100001F800600180060018006",
INIT_3D => X"00030C06600F0018000000001F8060018006001800600180060018006001F830",
INIT_3E => X"1FF87FE000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"C1FE06000C101FC00000000000000000000000000000000000038003001C0070"
)
	port map(
		SSR => '0',
		DI => "0",
		EN => '1',
		WE => '0',
		CLK => clk_i,
		ADDR => rom_addr_s(13 downto 0),
		DO => data0_s
	);

rom1: RAMB16_S1
	generic map(
INIT_00 => X"00000000003D830E1818606181860E0CD81E6001800600000001BE078C1C1860",
INIT_01 => X"60618186061C306F01800600000000003C030C081800600182060C300F000000",
INIT_02 => X"078000000000FC060C00180061FF860618301F00000000000000019E06CC1C18",
INIT_03 => X"3070618186061C306F0000000000000000180060018006001803F80180060030",
INIT_04 => X"180060000000018186061818606181860E0CD81E6001800607F030618006781B",
INIT_05 => X"0180060018006001F00000180060000000001800600180060018006001F00000",
INIT_06 => X"0018007C00000001818386039803E03983861818006001800600780300180060",
INIT_07 => X"66199866619986661BB83BA00000000000000018006001800600180060018006",
INIT_08 => X"0F00000000000000018186061818606181860E0CD81E60000000000000019986",
INIT_09 => X"830E1818606181860E0CD81E60000000000000003C030C181860618186060C30",
INIT_0A => X"D83E60000000180060019E06CC1C1860618186061C306F00000000001800603D",
INIT_0B => X"7F060618003C000F00060C181FC0000000000000000180060018006001860E18",
INIT_0C => X"1818606000000000000001E000C00180060018006001803F8018004000000000",
INIT_0D => X"001800F006601980C3030C18186060000000000000019E06CC1C186061818606",
INIT_0E => X"980C306060000000000000006601980FF036C199866618186060000000000000",
INIT_0F => X"30618006781B307061818606181860600000000000000181830C06600F003C01",
INIT_10 => X"03C00C003003C00E0000000001FF001800C006003001800C007FC000000007F0",
INIT_11 => X"800600180060018006001800600180060018006000000003800F000C003000F0",
INIT_12 => X"0000000F106EC11E0000000000000E007801800600F003C0018006001E003801",
INIT_13 => X"000000006003001800C007FE1FF830006000C001800000000000000000000000",
INIT_14 => X"404101040220070000000000000F007E01E807200F001800F001800600000000",
INIT_15 => X"0000001F8018006007E03FC08102F400000000000000000007003E0070022010",
INIT_16 => X"6F217883DE007800C0030000000036C1E7836C03C036C06600C0000000000000",
INIT_17 => X"000000000F807F018C0C183160C9838E07F01FC03E000000001F80C2052E1428",
INIT_18 => X"645FF0DB46DA06D00000000000000021008201B003004F217302E00240090018",
INIT_19 => X"000000000000800700F801800F006003000800600100000000001FF0BB45ED0A",
INIT_1A => X"17C859E1EB06BC0CE00F800C00000000000008005002E017C03E000000000000",
INIT_1B => X"D3FFCFFF00005002A00540050008005D80C900D8000000000000001C008C02CC",
INIT_1C => X"0000000600180000000000000000003FFC801200C9FD242C90D242C90D27ECBF",
INIT_1D => X"00000000000000000003001C00A007002801400E001000000000000000000000",
INIT_1E => X"86A619582AA11500A219186A619586AE0000000000007002600B803E00700000",
INIT_1F => X"FC3572A9C1FC00005552AA85552AA8555238CBEF0E38555071C71C11502A2191",
INIT_20 => X"AA85552AA800015542AB2FFC3572A9C1FC11502A219186061AB800015542AB2F",
INIT_21 => X"003800A001800000000000000000000000000000000FF05561FF800000005552",
INIT_22 => X"01FF87B413F85FE17F87B41FF83FC00000000000006003800A003800A003800A",
INIT_23 => X"EA1554AAA1554AAA0444444044444405C4494064446404444440444444000000",
INIT_24 => X"04001B013C07E007C07D83D00F6018000000001554AAA1554AAA15D4A9A1654A",
INIT_25 => X"07C01F000001C00700000008006003F01F601BC07F01A4038007000000000000",
INIT_26 => X"0000000000F8063010406300F800000000000000000057C0BF05000FC05F0080",
INIT_27 => X"FF00000FF06F60FF00000E7073819C84E6073839C00E0072001800E000000000",
INIT_28 => X"00000F807F018C0C183DE0C183DE04101DC03E00000FF06F60FF00000FF06F60",
INIT_29 => X"008087271FFC252000000000001F0086007003004C513C86761F6839C0420000",
INIT_2A => X"38044015405501FC17F03F800E80BA01B001000E001000000000000000000000",
INIT_2B => X"17A052814A07380FC02B00780E00618366CDFF1FAC3D607B0039019807C01D00",
INIT_2C => X"0040000073813B06E41EE033007F03B21CC86740E6000007780DC016015A05E8",
INIT_2D => X"CCCF33FFC7FE02401F805A00F000001B006C01500BA03F8028011007C00E0010",
INIT_2E => X"C00180000000006000C001800307FE1FF800C006003001801EF01B01AD86F633",
INIT_2F => X"13F07B011E04FC11A007800C0000000000006003001800C007FE1FF830006000",
INIT_30 => X"801E0000070013805801C007481E403E00E000B007C01A003804603BE1FC8278",
INIT_31 => X"FC0F7003C00F0024006003C006000007700D8036815A05E81FE03F007805400F",
INIT_32 => X"07000000001EF00F01BD86F612486FE1FF008807F01240FF8070020030018E07",
INIT_33 => X"83F70FDC11F03BC1F50B6024807C00000000780160073C0D581AA05581AC03E0",
INIT_34 => X"E863E0070000000007007E03BA09F8D7C1CA036C09B005400E0000182033004C",
INIT_35 => X"EC01A00F607541BB071C0C703F805701F000000E007C03B81CE0675198836E0D",
INIT_36 => X"045055206C00E0031C0EE01B006D01BC37D1D54D5717FC15503F807C04601980",
INIT_37 => X"631C81FA05EC1BB05D80C803200E401F00000C603B00FC03FE0FC83FA0FF03FE",
INIT_38 => X"EE07F00D401E00000DB03FC08101DC07702040AD03BC00103FC0DB000007807B",
INIT_39 => X"31C04201D011C46730FF81DC0080070008000000003DE03606FB1BEC4C91AEC3",
INIT_3A => X"C7771554777088800000000000C3056A0AD011814A851A14A81F800000000000",
INIT_3B => X"001FF0BB45ED0A645FF09985FF0DB46DA06D000000002221DDC5551DDC7771DD",
INIT_3C => X"0000000000000000000000000D806301DC0E383760DD838E077018C036000000",
INIT_3D => X"000005002B015E09E817E0BD81E407F00F0000000000007FE08302541EB83FC0",
INIT_3E => X"E0F301FA0BF006000000000000158054855E0B700E00DD038800000000000000",
INIT_3F => X"0000001E00C4062018007901FE03F000D802C00C0000001010011A80F00BF07C")
	port map(
		SSR => '0',
		DI => "0",
		EN => '1',
		WE => '0',
		CLK => clk_i,
		ADDR => rom_addr_s(13 downto 0),
		DO => data1_s);

rom2: RAMB16_S1
	generic map(
		INIT_00 => X"1BA06A81BA07180FC01E000000000300CB02280BA03FB07DC60E306801200000",
INIT_01 => X"C00000001CE0C606F71FBC3FF0FD441B10444000C00000000000000000780310",
INIT_02 => X"D01DC01400A803E0070008000003600F609783AC05C00F802A00A807F038E1C1",
INIT_03 => X"F01F800000C18306183060C3F607D800C00300180060030000000D8036007005",
INIT_04 => X"05D01FC036007002A00F80220000003000C00600181FC07F03180C6063018C07",
INIT_05 => X"001C000000002E609B027408E82EE0EE027C14E0210004000000000D80140174",
INIT_06 => X"D402D83EE0F587DC0070038006000000001DC03600D80BE837607F00F801C007",
INIT_07 => X"0FC03501FE00006300D803E00F801E008C05DA0AB01CC006003000007F00FA01",
INIT_08 => X"C3EB1FAC7EE0FA8BF0170000000000000000000004001000C003000E007801E0",
INIT_09 => X"80000000000000001800CC06A61BFC7FE1FA83DE00480000000000006031A0DD",
INIT_0A => X"FE01500000000000000000000000000000000008819281DE19F01F80F9019000",
INIT_0B => X"09C81E400000000000110055015407F05FC0FE003600F803C00600003FF864C0",
INIT_0C => X"007803F01DE067803F00B401E007800C0000000013C09C82D80EB037606B80DA",
INIT_0D => X"F807E036C0180000000000803B00B80BF817A1BF83E01E607600000000000000",
INIT_0E => X"18C07E00F30DFC3561E8067A0D780EC01000000000000018036C07E01F81FF81",
INIT_0F => X"83FE07F00F8000000000000F807F01240E383DE0F7830606301DC03E00000F78",
INIT_10 => X"000F807301940E183CE0FF83CE07F01CC03E000000006D30DD83FE0D28252094",
INIT_11 => X"02801C01BC1A418A88D101E01FE0C0C203081C11E27E0E40008003001C03C000",
INIT_12 => X"00000000000000000000000000000000000000000000040020008004001400A0",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"F860618186061818606000000000000000000000000000000000000000000000",
INIT_1C => X"000000000000000000000000000000000000000000000000000000600180FE0F",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0007FE1FF86060C3030C066019803C0060000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000")
	port map(
		SSR => '0',
		DI => "0",
		EN => '1',
		WE => '0',
		CLK => clk_i,
		ADDR => rom_addr_s(13 downto 0),
		DO => data2_s);

rom_addr_s <= std_logic_vector(to_unsigned(addr_i, rom_addr_s'length));
data_o <= data2_s when rom_addr_s(15 downto 14) = "10" else
	  data1_s when rom_addr_s(15 downto 14) = "01" else
	  data0_s;
end rtl;
